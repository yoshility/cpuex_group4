`default_nettype wire
module finv (
	input wire [31:0]  x,
  output wire [31:0] y,
  //output wire        ovf,
  input wire       clk,
  input wire       rstn
);
	wire      	sign = x[31];
	wire [ 7:0] exp_x = x[30:23];
	wire [22:0] frac_x = x[22:0];

	wire [ 9:0] addr = x[22:13];
	wire [12:0] dx = x[12:0];
	wire [35:0] dout;
	finv_table finv_table1(addr, dout, clk, rstn);

	wire [22:0] constant = dout[35:13];
	wire [12:0] gradient = dout[12:0];
	wire [25:0] dy_calc = gradient * dx;
	wire [22:0] frac_y = constant - dy_calc[25:3];

	wire [ 7:0] exp_x_unbiased = exp_x - 8'd127;
	wire [ 7:0] exp_y_unbiased = ~exp_x_unbiased + 8'd1;
	wire [ 7:0] exp_y = exp_y_unbiased + 8'd127;

	assign y = {sign , exp_y, frac_y};
endmodule

module fdiv (
	input  [31:0] x1,
	input  [31:0] x2,
	output [31:0] y,
	input 				clk,
	input					rstn
);
	wire [31:0] inv_x2;
	finv finv_in_fdiv(x2,inv_x2,clk,rstn);
	fmul fmul_in_fdiv(x1,inv_x2,y,clk,rstn);
endmodule

module finv_table (
	input		wire [ 9:0]	addr,
	output	reg  [35:0] dout,
	input 	wire 				clk,
	input 	wire 				rstn
);
	(*ram_style = "BLOCK"*) logic [35:0] finv_table [1023:0];
	always @(posedge clk) begin
		dout <= finv_table[addr];
	end
	initial begin
		finv_table[   0] = 36'b111111111011111111111111111111111000;
		finv_table[   1] = 36'b111111110011111111011111111111101000;
		finv_table[   2] = 36'b111111101011111110011111111111011000;
		finv_table[   3] = 36'b111111100100001101000011111111001000;
		finv_table[   4] = 36'b111111011100001011000001111110111000;
		finv_table[   5] = 36'b111111010100001000100011111110101000;
		finv_table[   6] = 36'b111111001100010101101001111110011001;
		finv_table[   7] = 36'b111111000100100010001111111110001001;
		finv_table[   8] = 36'b111110111100011110001111111101111001;
		finv_table[   9] = 36'b111110110100101001111001111101101010;
		finv_table[  10] = 36'b111110101101000101001101111101011011;
		finv_table[  11] = 36'b111110100100111111101101111101001011;
		finv_table[  12] = 36'b111110011101001001111001111100111011;
		finv_table[  13] = 36'b111110010101010011100101111100101100;
		finv_table[  14] = 36'b111110001101101101000001111100011101;
		finv_table[  15] = 36'b111110000101110101101111111100001101;
		finv_table[  16] = 36'b111101111110001110001111111011111110;
		finv_table[  17] = 36'b111101110110010110000001111011101111;
		finv_table[  18] = 36'b111101101110011101010011111011011111;
		finv_table[  19] = 36'b111101100111000100101101111011010001;
		finv_table[  20] = 36'b111101011111001011000001111011000001;
		finv_table[  21] = 36'b111101010111100001001011111010110010;
		finv_table[  22] = 36'b111101001111110110110111111010100011;
		finv_table[  23] = 36'b111101001000001100000101111010010100;
		finv_table[  24] = 36'b111101000000100000110101111010000101;
		finv_table[  25] = 36'b111100111001000101011111111001110111;
		finv_table[  26] = 36'b111100110001011001010011111001101000;
		finv_table[  27] = 36'b111100101001101100101001111001011001;
		finv_table[  28] = 36'b111100100010001111111101111001001010;
		finv_table[  29] = 36'b111100011010100010010111111000111011;
		finv_table[  30] = 36'b111100010011000100110001111000101101;
		finv_table[  31] = 36'b111100001011010110001111111000011110;
		finv_table[  32] = 36'b111100000100001000001111111000010000;
		finv_table[  33] = 36'b111011111100011000110001111000000001;
		finv_table[  34] = 36'b111011110101001001111001110111110011;
		finv_table[  35] = 36'b111011101101011001011111110111100100;
		finv_table[  36] = 36'b111011100110001001101111110111010110;
		finv_table[  37] = 36'b111011011110101000111101110111000111;
		finv_table[  38] = 36'b111011010111000111110001110110111001;
		finv_table[  39] = 36'b111011001111100110000101110110101010;
		finv_table[  40] = 36'b111011001000010100100101110110011100;
		finv_table[  41] = 36'b111011000001000010101001110110001110;
		finv_table[  42] = 36'b111010111001011111100111110110000000;
		finv_table[  43] = 36'b111010110010001100110011110101110010;
		finv_table[  44] = 36'b111010101010111001100011110101100100;
		finv_table[  45] = 36'b111010100011010101001001110101010101;
		finv_table[  46] = 36'b111010011100010001110001110101001000;
		finv_table[  47] = 36'b111010010100111101001101110100111010;
		finv_table[  48] = 36'b111010001101010111011101110100101011;
		finv_table[  49] = 36'b111010000110010010110001110100011110;
		finv_table[  50] = 36'b111001111110111100111001110100010000;
		finv_table[  51] = 36'b111001110111110111011001110100000010;
		finv_table[  52] = 36'b111001110000100000100111110011110100;
		finv_table[  53] = 36'b111001101001001001011101110011100110;
		finv_table[  54] = 36'b111001100010000010101001110011011001;
		finv_table[  55] = 36'b111001011010111011011101110011001011;
		finv_table[  56] = 36'b111001010011100010111101110010111101;
		finv_table[  57] = 36'b111001001100011010111001110010110000;
		finv_table[  58] = 36'b111001000101010010011011110010100010;
		finv_table[  59] = 36'b111000111110001001100011110010010101;
		finv_table[  60] = 36'b111000110111000000001111110010000111;
		finv_table[  61] = 36'b111000101111110110100001110001111010;
		finv_table[  62] = 36'b111000101000111101010101110001101101;
		finv_table[  63] = 36'b111000100001100001110001110001011111;
		finv_table[  64] = 36'b111000011010100111110001110001010010;
		finv_table[  65] = 36'b111000010011011100010101110001000100;
		finv_table[  66] = 36'b111000001100100001100001110000110111;
		finv_table[  67] = 36'b111000000101010101010001110000101010;
		finv_table[  68] = 36'b110111111110011001101001110000011101;
		finv_table[  69] = 36'b110111110111001100100001110000001111;
		finv_table[  70] = 36'b110111110000100001001101110000000011;
		finv_table[  71] = 36'b110111101001010011001101101111110101;
		finv_table[  72] = 36'b110111100010010101111101101111101000;
		finv_table[  73] = 36'b110111011011011000010011101111011011;
		finv_table[  74] = 36'b110111010100011010001111101111001110;
		finv_table[  75] = 36'b110111001101011011110001101111000001;
		finv_table[  76] = 36'b110111000110011100111001101110110100;
		finv_table[  77] = 36'b110110111111101110110101101110101000;
		finv_table[  78] = 36'b110110111000101111001001101110011011;
		finv_table[  79] = 36'b110110110001101111000011101110001110;
		finv_table[  80] = 36'b110110101010111111110011101110000001;
		finv_table[  81] = 36'b110110100011111110111001101101110100;
		finv_table[  82] = 36'b110110011101001110110111101101101000;
		finv_table[  83] = 36'b110110010110011110011011101101011011;
		finv_table[  84] = 36'b110110001111011100010011101101001110;
		finv_table[  85] = 36'b110110001000101011000111101101000010;
		finv_table[  86] = 36'b110110000001111001100001101100110101;
		finv_table[  87] = 36'b110101111011000111100001101100101001;
		finv_table[  88] = 36'b110101110100010101001001101100011100;
		finv_table[  89] = 36'b110101101101100010011001101100010000;
		finv_table[  90] = 36'b110101100111000000101001101100000100;
		finv_table[  91] = 36'b110101011111111011101101101011110111;
		finv_table[  92] = 36'b110101011001011001001101101011101011;
		finv_table[  93] = 36'b110101010010100100110111101011011110;
		finv_table[  94] = 36'b110101001011110000001001101011010010;
		finv_table[  95] = 36'b110101000101001100100001101011000110;
		finv_table[  96] = 36'b110100111110101000100001101010111010;
		finv_table[  97] = 36'b110100110111110010100111101010101101;
		finv_table[  98] = 36'b110100110000111100010101101010100001;
		finv_table[  99] = 36'b110100101010101000101111101010010101;
		finv_table[ 100] = 36'b110100100011110001101101101010001001;
		finv_table[ 101] = 36'b110100011101001011110101101001111101;
		finv_table[ 102] = 36'b110100010110100101100101101001110001;
		finv_table[ 103] = 36'b110100010000010000100011101001100101;
		finv_table[ 104] = 36'b110100001001010111111101101001011001;
		finv_table[ 105] = 36'b110100000010110000100101101001001101;
		finv_table[ 106] = 36'b110011111100001000110101101001000001;
		finv_table[ 107] = 36'b110011110101110010010101101000110101;
		finv_table[ 108] = 36'b110011101111001001110111101000101001;
		finv_table[ 109] = 36'b110011101000110010101011101000011110;
		finv_table[ 110] = 36'b110011100001110111101101101000010001;
		finv_table[ 111] = 36'b110011011011110001100101101000000110;
		finv_table[ 112] = 36'b110011010101000111100011100111111010;
		finv_table[ 113] = 36'b110011001110011101001101100111101110;
		finv_table[ 114] = 36'b110011001000000100001101100111100011;
		finv_table[ 115] = 36'b110011000001101010110111100111010111;
		finv_table[ 116] = 36'b110010111011010001001101100111001100;
		finv_table[ 117] = 36'b110010110100110111001001100111000000;
		finv_table[ 118] = 36'b110010101110001010111001100110110100;
		finv_table[ 119] = 36'b110010101000000001111111100110101001;
		finv_table[ 120] = 36'b110010100001010101000001100110011101;
		finv_table[ 121] = 36'b110010011011001011011001100110010010;
		finv_table[ 122] = 36'b110010010100101111100101100110000111;
		finv_table[ 123] = 36'b110010001110010011010101100101111011;
		finv_table[ 124] = 36'b110010001000001000101101100101110000;
		finv_table[ 125] = 36'b110010000001011001110111100101100100;
		finv_table[ 126] = 36'b110001111011001110100011100101011001;
		finv_table[ 127] = 36'b110001110101000010111001100101001110;
		finv_table[ 128] = 36'b110001101110100100111001100101000011;
		finv_table[ 129] = 36'b110001101000011000100011100100111000;
		finv_table[ 130] = 36'b110001100001111001110101100100101100;
		finv_table[ 131] = 36'b110001011011101100110001100100100001;
		finv_table[ 132] = 36'b110001010101011111011001100100010110;
		finv_table[ 133] = 36'b110001001111010001101101100100001011;
		finv_table[ 134] = 36'b110001001000110001100011100100000000;
		finv_table[ 135] = 36'b110001000010110101001111100011110101;
		finv_table[ 136] = 36'b110000111100010100010111100011101010;
		finv_table[ 137] = 36'b110000110110010111011001100011011111;
		finv_table[ 138] = 36'b110000101111110101110101100011010100;
		finv_table[ 139] = 36'b110000101001111000001101100011001001;
		finv_table[ 140] = 36'b110000100011101000000101100010111110;
		finv_table[ 141] = 36'b110000011101010111100111100010110011;
		finv_table[ 142] = 36'b110000010111011001000001100010101001;
		finv_table[ 143] = 36'b110000010001000111110111100010011110;
		finv_table[ 144] = 36'b110000001010110110011001100010010011;
		finv_table[ 145] = 36'b110000000100110110110011100010001000;
		finv_table[ 146] = 36'b101111111110110110111001100001111110;
		finv_table[ 147] = 36'b101111111000100100010111100001110011;
		finv_table[ 148] = 36'b101111110010010001011111100001101000;
		finv_table[ 149] = 36'b101111101100100010111011100001011110;
		finv_table[ 150] = 36'b101111100110001111010111100001010011;
		finv_table[ 151] = 36'b101111100000001101110101100001001000;
		finv_table[ 152] = 36'b101111011010001011111101100000111110;
		finv_table[ 153] = 36'b101111010011110111010101100000110011;
		finv_table[ 154] = 36'b101111001110000111001101100000101001;
		finv_table[ 155] = 36'b101111001000000100010111100000011110;
		finv_table[ 156] = 36'b101111000010000001001011100000010100;
		finv_table[ 157] = 36'b101110111011111101101001100000001001;
		finv_table[ 158] = 36'b101110110101111001110101011111111111;
		finv_table[ 159] = 36'b101110101111110101101001011111110100;
		finv_table[ 160] = 36'b101110101010000011101001011111101010;
		finv_table[ 161] = 36'b101110100011111110110011011111100000;
		finv_table[ 162] = 36'b101110011110001100001011011111010110;
		finv_table[ 163] = 36'b101110011000000110101101011111001011;
		finv_table[ 164] = 36'b101110010010000000111001011111000001;
		finv_table[ 165] = 36'b101110001100001101010101011110110111;
		finv_table[ 166] = 36'b101110000110011001011101011110101101;
		finv_table[ 167] = 36'b101110000000010010101001011110100010;
		finv_table[ 168] = 36'b101101111010011110001001011110011000;
		finv_table[ 169] = 36'b101101110100101001010101011110001110;
		finv_table[ 170] = 36'b101101101110100001100011011110000100;
		finv_table[ 171] = 36'b101101101000111110110011011101111010;
		finv_table[ 172] = 36'b101101100010110110010111011101110000;
		finv_table[ 173] = 36'b101101011101010011000001011101100110;
		finv_table[ 174] = 36'b101101010111001001111001011101011100;
		finv_table[ 175] = 36'b101101010001010011001101011101010010;
		finv_table[ 176] = 36'b101101001011101110111101011101001000;
		finv_table[ 177] = 36'b101101000101110111101001011100111110;
		finv_table[ 178] = 36'b101100111111101101010001011100110100;
		finv_table[ 179] = 36'b101100111010011010111001011100101011;
		finv_table[ 180] = 36'b101100110100001111110101011100100000;
		finv_table[ 181] = 36'b101100101110101010000101011100010111;
		finv_table[ 182] = 36'b101100101000110001001101011100001101;
		finv_table[ 183] = 36'b101100100011001010111001011100000011;
		finv_table[ 184] = 36'b101100011101010001011001011011111001;
		finv_table[ 185] = 36'b101100010111101010011111011011110000;
		finv_table[ 186] = 36'b101100010001110000010111011011100110;
		finv_table[ 187] = 36'b101100001100001000110101011011011100;
		finv_table[ 188] = 36'b101100000110100001000001011011010011;
		finv_table[ 189] = 36'b101100000000111000111001011011001001;
		finv_table[ 190] = 36'b101011111010111101100011011010111111;
		finv_table[ 191] = 36'b101011110101010100110101011010110110;
		finv_table[ 192] = 36'b101011101111101011110101011010101100;
		finv_table[ 193] = 36'b101011101010000010100011011010100011;
		finv_table[ 194] = 36'b101011100100011000111101011010011001;
		finv_table[ 195] = 36'b101011011110101111000101011010010000;
		finv_table[ 196] = 36'b101011011001000100110111011010000110;
		finv_table[ 197] = 36'b101011010011011010011001011001111101;
		finv_table[ 198] = 36'b101011001110000010101101011001110100;
		finv_table[ 199] = 36'b101011001000000100100001011001101010;
		finv_table[ 200] = 36'b101011000010101100010001011001100001;
		finv_table[ 201] = 36'b101010111101000000100101011001010111;
		finv_table[ 202] = 36'b101010110111100111110001011001001110;
		finv_table[ 203] = 36'b101010110001111011100001011001000101;
		finv_table[ 204] = 36'b101010101100001110111101011000111011;
		finv_table[ 205] = 36'b101010100110110101010011011000110010;
		finv_table[ 206] = 36'b101010100001001000001001011000101001;
		finv_table[ 207] = 36'b101010011011101101111011011000100000;
		finv_table[ 208] = 36'b101010010110010011011011011000010111;
		finv_table[ 209] = 36'b101010010000100101011001011000001101;
		finv_table[ 210] = 36'b101010001011001010010011011000000100;
		finv_table[ 211] = 36'b101010000101011011101011010111111011;
		finv_table[ 212] = 36'b101010000000010011010101010111110010;
		finv_table[ 213] = 36'b101001111010100100001001010111101001;
		finv_table[ 214] = 36'b101001110101011011010001010111100000;
		finv_table[ 215] = 36'b101001101111101011011101010111010111;
		finv_table[ 216] = 36'b101001101010001110101101010111001110;
		finv_table[ 217] = 36'b101001100100110001101011010111000101;
		finv_table[ 218] = 36'b101001011111010100010111010110111100;
		finv_table[ 219] = 36'b101001011010001010001011010110110011;
		finv_table[ 220] = 36'b101001010100011000111001010110101010;
		finv_table[ 221] = 36'b101001001111001110001001010110100001;
		finv_table[ 222] = 36'b101001001001101111101101010110011000;
		finv_table[ 223] = 36'b101001000100010001000001010110001111;
		finv_table[ 224] = 36'b101000111111000101100001010110000111;
		finv_table[ 225] = 36'b101000111001100110001111010101111110;
		finv_table[ 226] = 36'b101000110100000110101011010101110101;
		finv_table[ 227] = 36'b101000101110111010011001010101101100;
		finv_table[ 228] = 36'b101000101001011010010001010101100011;
		finv_table[ 229] = 36'b101000100100001101011011010101011011;
		finv_table[ 230] = 36'b101000011110101100101111010101010010;
		finv_table[ 231] = 36'b101000011001011111010111010101001001;
		finv_table[ 232] = 36'b101000010100010001110001010101000001;
		finv_table[ 233] = 36'b101000001110110000001101010100111000;
		finv_table[ 234] = 36'b101000001001100010000101010100101111;
		finv_table[ 235] = 36'b101000000100010011101001010100100111;
		finv_table[ 236] = 36'b100111111111000100111101010100011110;
		finv_table[ 237] = 36'b100111111001100010010001010100010101;
		finv_table[ 238] = 36'b100111110100100110110011010100001101;
		finv_table[ 239] = 36'b100111101111000011100101010100000100;
		finv_table[ 240] = 36'b100111101010000111100101010011111100;
		finv_table[ 241] = 36'b100111100100100011110001010011110011;
		finv_table[ 242] = 36'b100111011111100111010011010011101011;
		finv_table[ 243] = 36'b100111011010000010111101010011100010;
		finv_table[ 244] = 36'b100111010101000101111101010011011010;
		finv_table[ 245] = 36'b100111001111110100111001010011010010;
		finv_table[ 246] = 36'b100111001010100011100001010011001001;
		finv_table[ 247] = 36'b100111000101100101110001010011000001;
		finv_table[ 248] = 36'b100111000000000000000001010010111000;
		finv_table[ 249] = 36'b100110111011000001110001010010110000;
		finv_table[ 250] = 36'b100110110110000011010001010010101000;
		finv_table[ 251] = 36'b100110110000110000100111010010100000;
		finv_table[ 252] = 36'b100110101011011101101101010010010111;
		finv_table[ 253] = 36'b100110100110011110011011010010001111;
		finv_table[ 254] = 36'b100110100001001010111101010010000111;
		finv_table[ 255] = 36'b100110011100001011001101010001111111;
		finv_table[ 256] = 36'b100110010111001011001101010001110111;
		finv_table[ 257] = 36'b100110010001110110111101010001101110;
		finv_table[ 258] = 36'b100110001100110110011101010001100110;
		finv_table[ 259] = 36'b100110000111110101101101010001011110;
		finv_table[ 260] = 36'b100110000010100000101001010001010110;
		finv_table[ 261] = 36'b100101111101011111011001010001001110;
		finv_table[ 262] = 36'b100101111000011101111001010001000110;
		finv_table[ 263] = 36'b100101110011011100001001010000111110;
		finv_table[ 264] = 36'b100101101110011010001001010000110110;
		finv_table[ 265] = 36'b100101101001010111111001010000101110;
		finv_table[ 266] = 36'b100101100100010101011001010000100110;
		finv_table[ 267] = 36'b100101011111010010101001010000011110;
		finv_table[ 268] = 36'b100101011010001111101001010000010110;
		finv_table[ 269] = 36'b100101010101001100011001010000001110;
		finv_table[ 270] = 36'b100101010000001000111001010000000110;
		finv_table[ 271] = 36'b100101001011000101001001001111111110;
		finv_table[ 272] = 36'b100101000110010101011001001111110110;
		finv_table[ 273] = 36'b100101000000111100110111001111101110;
		finv_table[ 274] = 36'b100100111100100000111011001111100111;
		finv_table[ 275] = 36'b100100110111000111111001001111011110;
		finv_table[ 276] = 36'b100100110010010111001101001111010111;
		finv_table[ 277] = 36'b100100101101010001111101001111001111;
		finv_table[ 278] = 36'b100100101000100000110011001111000111;
		finv_table[ 279] = 36'b100100100011011011000001001110111111;
		finv_table[ 280] = 36'b100100011110010101000011001110110111;
		finv_table[ 281] = 36'b100100011001100011001011001110110000;
		finv_table[ 282] = 36'b100100010100110001000101001110101000;
		finv_table[ 283] = 36'b100100001111101010010101001110100000;
		finv_table[ 284] = 36'b100100001010110111110001001110011001;
		finv_table[ 285] = 36'b100100000110000100111101001110010001;
		finv_table[ 286] = 36'b100100000000111101011101001110001001;
		finv_table[ 287] = 36'b100011111100011110101101001110000010;
		finv_table[ 288] = 36'b100011110111000010001101001101111010;
		finv_table[ 289] = 36'b100011110010100010111101001101110011;
		finv_table[ 290] = 36'b100011101101101111000001001101101011;
		finv_table[ 291] = 36'b100011101000100110010001001101100011;
		finv_table[ 292] = 36'b100011100100000110011001001101011100;
		finv_table[ 293] = 36'b100011011110111101001001001101010100;
		finv_table[ 294] = 36'b100011011010001000001101001101001101;
		finv_table[ 295] = 36'b100011010101100111101101001101000110;
		finv_table[ 296] = 36'b100011010000011101101101001100111110;
		finv_table[ 297] = 36'b100011001011111100101101001100110111;
		finv_table[ 298] = 36'b100011000110110010001101001100101111;
		finv_table[ 299] = 36'b100011000010010000110101001100101000;
		finv_table[ 300] = 36'b100010111101011010100001001100100000;
		finv_table[ 301] = 36'b100010111000100011111101001100011001;
		finv_table[ 302] = 36'b100010110100000001111001001100010010;
		finv_table[ 303] = 36'b100010101111001010111001001100001010;
		finv_table[ 304] = 36'b100010101010010011101001001100000011;
		finv_table[ 305] = 36'b100010100101011100001001001011111011;
		finv_table[ 306] = 36'b100010100000111001001101001011110100;
		finv_table[ 307] = 36'b100010011100000001010001001011101101;
		finv_table[ 308] = 36'b100010010111011101111001001011100110;
		finv_table[ 309] = 36'b100010010010100101011101001011011110;
		finv_table[ 310] = 36'b100010001110000001101001001011010111;
		finv_table[ 311] = 36'b100010001001001000110001001011010000;
		finv_table[ 312] = 36'b100010000100100100100001001011001001;
		finv_table[ 313] = 36'b100010000000000000000001001011000010;
		finv_table[ 314] = 36'b100001111011000110011101001010111010;
		finv_table[ 315] = 36'b100001110110100001100001001010110011;
		finv_table[ 316] = 36'b100001110001111100011001001010101100;
		finv_table[ 317] = 36'b100001101101000010000111001010100101;
		finv_table[ 318] = 36'b100001101000011100100011001010011110;
		finv_table[ 319] = 36'b100001100011110110110001001010010111;
		finv_table[ 320] = 36'b100001011111010000110001001010010000;
		finv_table[ 321] = 36'b100001011010101010100011001010001001;
		finv_table[ 322] = 36'b100001010101101111000101001010000001;
		finv_table[ 323] = 36'b100001010001011101011101001001111011;
		finv_table[ 324] = 36'b100001001100100001100011001001110011;
		finv_table[ 325] = 36'b100001001000001111100001001001101101;
		finv_table[ 326] = 36'b100001000011101000001101001001100110;
		finv_table[ 327] = 36'b100000111110101011100101001001011110;
		finv_table[ 328] = 36'b100000111010011000111101001001011000;
		finv_table[ 329] = 36'b100000110101110000111101001001010001;
		finv_table[ 330] = 36'b100000110001001000110011001001001010;
		finv_table[ 331] = 36'b100000101100100000011001001001000011;
		finv_table[ 332] = 36'b100000100111110111110001001000111100;
		finv_table[ 333] = 36'b100000100011100100000111001000110101;
		finv_table[ 334] = 36'b100000011110111011000011001000101110;
		finv_table[ 335] = 36'b100000011010010001110001001000100111;
		finv_table[ 336] = 36'b100000010101111101100001001000100001;
		finv_table[ 337] = 36'b100000010001010011110011001000011010;
		finv_table[ 338] = 36'b100000001100101001110111001000010011;
		finv_table[ 339] = 36'b100000001000010101000001001000001100;
		finv_table[ 340] = 36'b100000000011101010101001001000000101;
		finv_table[ 341] = 36'b011111111111010101010111000111111111;
		finv_table[ 342] = 36'b011111111010101010100011000111111000;
		finv_table[ 343] = 36'b011111110110010100111001000111110001;
		finv_table[ 344] = 36'b011111110001101001101001000111101010;
		finv_table[ 345] = 36'b011111101101101000111101000111100100;
		finv_table[ 346] = 36'b011111101000100111110101000111011101;
		finv_table[ 347] = 36'b011111100100010001011001000111010110;
		finv_table[ 348] = 36'b011111011111111010101011000111010000;
		finv_table[ 349] = 36'b011111011011100011110001000111001001;
		finv_table[ 350] = 36'b011111010111001100101101000111000011;
		finv_table[ 351] = 36'b011111010010011111111011000110111100;
		finv_table[ 352] = 36'b011111001110001000011011000110110101;
		finv_table[ 353] = 36'b011111001001110000101101000110101111;
		finv_table[ 354] = 36'b011111000101011000110011000110101000;
		finv_table[ 355] = 36'b011111000000101011001001000110100001;
		finv_table[ 356] = 36'b011110111100101000011001000110011011;
		finv_table[ 357] = 36'b011110111000001111111001000110010101;
		finv_table[ 358] = 36'b011110110011100001100101000110001110;
		finv_table[ 359] = 36'b011110101111011110010001000110001000;
		finv_table[ 360] = 36'b011110101010101111100001000110000001;
		finv_table[ 361] = 36'b011110100110101011110101000101111011;
		finv_table[ 362] = 36'b011110100010010010010001000101110100;
		finv_table[ 363] = 36'b011110011101111000100011000101101110;
		finv_table[ 364] = 36'b011110011001011110101001000101100111;
		finv_table[ 365] = 36'b011110010101000100011101000101100001;
		finv_table[ 366] = 36'b011110010000101010001001000101011010;
		finv_table[ 367] = 36'b011110001100100101010101000101010100;
		finv_table[ 368] = 36'b011110001000001010100101000101001110;
		finv_table[ 369] = 36'b011110000011101111100111000101000111;
		finv_table[ 370] = 36'b011101111111101010010001000101000001;
		finv_table[ 371] = 36'b011101111010111001000101000100111010;
		finv_table[ 372] = 36'b011101110111001001001001000100110101;
		finv_table[ 373] = 36'b011101110010010111100011000100101110;
		finv_table[ 374] = 36'b011101101110010001011011000100101000;
		finv_table[ 375] = 36'b011101101010001011000111000100100010;
		finv_table[ 376] = 36'b011101100101101110110001000100011011;
		finv_table[ 377] = 36'b011101100001010010001001000100010101;
		finv_table[ 378] = 36'b011101011101001011010001000100001111;
		finv_table[ 379] = 36'b011101011001000100001101000100001001;
		finv_table[ 380] = 36'b011101010100100111000001000100000010;
		finv_table[ 381] = 36'b011101010000011111100111000011111100;
		finv_table[ 382] = 36'b011101001100000010000001000011110110;
		finv_table[ 383] = 36'b011101000111111010001101000011110000;
		finv_table[ 384] = 36'b011101000011110010001101000011101010;
		finv_table[ 385] = 36'b011100111111101010000001000011100100;
		finv_table[ 386] = 36'b011100111011001011100111000011011101;
		finv_table[ 387] = 36'b011100110111000011000001000011010111;
		finv_table[ 388] = 36'b011100110010111010010011000011010001;
		finv_table[ 389] = 36'b011100101110011011010001000011001011;
		finv_table[ 390] = 36'b011100101010101000010001000011000101;
		finv_table[ 391] = 36'b011100100110001000110101000010111111;
		finv_table[ 392] = 36'b011100100001111111010101000010111001;
		finv_table[ 393] = 36'b011100011101110101101001000010110011;
		finv_table[ 394] = 36'b011100011010000001111011000010101101;
		finv_table[ 395] = 36'b011100010101100001101101000010100111;
		finv_table[ 396] = 36'b011100010001010111011101000010100001;
		finv_table[ 397] = 36'b011100001101001101000001000010011011;
		finv_table[ 398] = 36'b011100001001000010011001000010010101;
		finv_table[ 399] = 36'b011100000100110111100101000010001111;
		finv_table[ 400] = 36'b011100000000101100100011000010001001;
		finv_table[ 401] = 36'b011011111100110111101001000010000011;
		finv_table[ 402] = 36'b011011111000101100010001000001111101;
		finv_table[ 403] = 36'b011011110100001010011001000001110111;
		finv_table[ 404] = 36'b011011110000010100111101000001110001;
		finv_table[ 405] = 36'b011011101100001001000001000001101011;
		finv_table[ 406] = 36'b011011101000010011001111000001100110;
		finv_table[ 407] = 36'b011011100100000110111011000001100000;
		finv_table[ 408] = 36'b011011011111111010011011000001011010;
		finv_table[ 409] = 36'b011011011011101101101111000001010100;
		finv_table[ 410] = 36'b011011010111110111010001000001001110;
		finv_table[ 411] = 36'b011011010011101010001101000001001000;
		finv_table[ 412] = 36'b011011001111011100111101000001000010;
		finv_table[ 413] = 36'b011011001011100101111101000000111101;
		finv_table[ 414] = 36'b011011000111011000010101000000110111;
		finv_table[ 415] = 36'b011011000011100001000001000000110001;
		finv_table[ 416] = 36'b011010111111101001100001000000101100;
		finv_table[ 417] = 36'b011010111011000100110101000000100101;
		finv_table[ 418] = 36'b011010110111100011100001000000100000;
		finv_table[ 419] = 36'b011010110011010100111101000000011010;
		finv_table[ 420] = 36'b011010101111000110001101000000010100;
		finv_table[ 421] = 36'b011010101011001101110101000000001111;
		finv_table[ 422] = 36'b011010100111010101010101000000001001;
		finv_table[ 423] = 36'b011010100011000101111111000000000011;
		finv_table[ 424] = 36'b011010011111100011101110111111111110;
		finv_table[ 425] = 36'b011010011010111101011010111111111000;
		finv_table[ 426] = 36'b011010010111011010110100111111110011;
		finv_table[ 427] = 36'b011010010011001010110000111111101101;
		finv_table[ 428] = 36'b011010001111010001001110111111100111;
		finv_table[ 429] = 36'b011010001011010111011110111111100010;
		finv_table[ 430] = 36'b011010000111011101100100111111011100;
		finv_table[ 431] = 36'b011010000011001100110000111111010110;
		finv_table[ 432] = 36'b011001111111101001010000111111010001;
		finv_table[ 433] = 36'b011001111011011000000100111111001011;
		finv_table[ 434] = 36'b011001110111011101011110111111000110;
		finv_table[ 435] = 36'b011001110011100010101110111111000000;
		finv_table[ 436] = 36'b011001101111100111110000111110111011;
		finv_table[ 437] = 36'b011001101011101100101010111110110101;
		finv_table[ 438] = 36'b011001101000001000001110111110110000;
		finv_table[ 439] = 36'b011001100011110101111100111110101010;
		finv_table[ 440] = 36'b011001011111111010010100111110100101;
		finv_table[ 441] = 36'b011001011011111110100000111110011111;
		finv_table[ 442] = 36'b011001011000000010100000111110011010;
		finv_table[ 443] = 36'b011001010100011101010100111110010101;
		finv_table[ 444] = 36'b011001010000001010000100111110001111;
		finv_table[ 445] = 36'b011001001100100100100000111110001010;
		finv_table[ 446] = 36'b011001001000100111111000111110000100;
		finv_table[ 447] = 36'b011001000100101011000100111101111111;
		finv_table[ 448] = 36'b011001000001000101000010111101111010;
		finv_table[ 449] = 36'b011000111100110000110110111101110100;
		finv_table[ 450] = 36'b011000111001001010100100111101101111;
		finv_table[ 451] = 36'b011000110101001101000000111101101001;
		finv_table[ 452] = 36'b011000110001100110011000111101100100;
		finv_table[ 453] = 36'b011000101101101000100100111101011111;
		finv_table[ 454] = 36'b011000101001101010100010111101011001;
		finv_table[ 455] = 36'b011000100101101100010100111101010100;
		finv_table[ 456] = 36'b011000100010000101000100111101001111;
		finv_table[ 457] = 36'b011000011110011101101010111101001010;
		finv_table[ 458] = 36'b011000011010000111110010111101000100;
		finv_table[ 459] = 36'b011000010110110111001110111100111111;
		finv_table[ 460] = 36'b011000010010111000001010111100111010;
		finv_table[ 461] = 36'b011000001110111000111100111100110100;
		finv_table[ 462] = 36'b011000001011010000110000111100101111;
		finv_table[ 463] = 36'b011000000111010001001010111100101010;
		finv_table[ 464] = 36'b011000000011101000101100111100100101;
		finv_table[ 465] = 36'b010111111111101000110000111100011111;
		finv_table[ 466] = 36'b010111111100010111001100111100011011;
		finv_table[ 467] = 36'b010111110111111111101000111100010101;
		finv_table[ 468] = 36'b010111110100101101110100111100010000;
		finv_table[ 469] = 36'b010111110000101101010000111100001011;
		finv_table[ 470] = 36'b010111101101000011110010111100000110;
		finv_table[ 471] = 36'b010111101001000010110110111100000000;
		finv_table[ 472] = 36'b010111100101011001000110111011111011;
		finv_table[ 473] = 36'b010111100001101111001100111011110110;
		finv_table[ 474] = 36'b010111011110000101001000111011110001;
		finv_table[ 475] = 36'b010111011010011010111010111011101100;
		finv_table[ 476] = 36'b010111010110011001000100111011100111;
		finv_table[ 477] = 36'b010111010011000110000000111011100010;
		finv_table[ 478] = 36'b010111001111000011111000111011011101;
		finv_table[ 479] = 36'b010111001011011001000000111011011000;
		finv_table[ 480] = 36'b010111000111101110000000111011010011;
		finv_table[ 481] = 36'b010111000011101011010100111011001101;
		finv_table[ 482] = 36'b010111000000010111100100111011001001;
		finv_table[ 483] = 36'b010110111100101100000110111011000100;
		finv_table[ 484] = 36'b010110111000101000111000111010111110;
		finv_table[ 485] = 36'b010110110101010100101100111010111010;
		finv_table[ 486] = 36'b010110110001101000110000111010110101;
		finv_table[ 487] = 36'b010110101101111100101010111010110000;
		finv_table[ 488] = 36'b010110101001111000110010111010101010;
		finv_table[ 489] = 36'b010110100110100100000000111010100110;
		finv_table[ 490] = 36'b010110100010110111011100111010100001;
		finv_table[ 491] = 36'b010110011111001010110000111010011100;
		finv_table[ 492] = 36'b010110011011110101100100111010010111;
		finv_table[ 493] = 36'b010110010111110000110100111010010010;
		finv_table[ 494] = 36'b010110010100011011011000111010001101;
		finv_table[ 495] = 36'b010110010000010110010010111010001000;
		finv_table[ 496] = 36'b010110001101000000100010111010000011;
		finv_table[ 497] = 36'b010110001001101010101000111001111111;
		finv_table[ 498] = 36'b010110000101100101000100111001111001;
		finv_table[ 499] = 36'b010110000010001110111000111001110101;
		finv_table[ 500] = 36'b010101111110100000110000111001110000;
		finv_table[ 501] = 36'b010101111010110010011100111001101011;
		finv_table[ 502] = 36'b010101110111011011111000111001100110;
		finv_table[ 503] = 36'b010101110011101101010000111001100001;
		finv_table[ 504] = 36'b010101110000010110011000111001011101;
		finv_table[ 505] = 36'b010101101100001111100110111001010111;
		finv_table[ 506] = 36'b010101101001010000011000111001010011;
		finv_table[ 507] = 36'b010101100101001001001110111001001110;
		finv_table[ 508] = 36'b010101100001110001110010111001001001;
		finv_table[ 509] = 36'b010101011110011010001100111001000101;
		finv_table[ 510] = 36'b010101011010101010100000111001000000;
		finv_table[ 511] = 36'b010101010110111010101100111000111011;
		finv_table[ 512] = 36'b010101010011100010101010111000110110;
		finv_table[ 513] = 36'b010101010000001010100010111000110010;
		finv_table[ 514] = 36'b010101001100011010001100111000101101;
		finv_table[ 515] = 36'b010101001001000001110100111000101000;
		finv_table[ 516] = 36'b010101000101010001001100111000100011;
		finv_table[ 517] = 36'b010101000001111000011100111000011111;
		finv_table[ 518] = 36'b010100111110011111101000111000011010;
		finv_table[ 519] = 36'b010100111010101110100010111000010101;
		finv_table[ 520] = 36'b010100110111010101011000111000010001;
		finv_table[ 521] = 36'b010100110011100100000000111000001100;
		finv_table[ 522] = 36'b010100110000001010100110111000000111;
		finv_table[ 523] = 36'b010100101100110001000100111000000011;
		finv_table[ 524] = 36'b010100101001010111010110110111111110;
		finv_table[ 525] = 36'b010100100101100101010100110111111001;
		finv_table[ 526] = 36'b010100100010100011100100110111110101;
		finv_table[ 527] = 36'b010100011110110001010000110111110000;
		finv_table[ 528] = 36'b010100011010111110110000110111101011;
		finv_table[ 529] = 36'b010100010111111100100110110111100111;
		finv_table[ 530] = 36'b010100010100100010000100110111100011;
		finv_table[ 531] = 36'b010100010000101111000110110111011110;
		finv_table[ 532] = 36'b010100001101010100010100110111011001;
		finv_table[ 533] = 36'b010100001001111001010100110111010101;
		finv_table[ 534] = 36'b010100000110011110010000110111010000;
		finv_table[ 535] = 36'b010100000011000011000000110111001100;
		finv_table[ 536] = 36'b010011111111100111101000110111000111;
		finv_table[ 537] = 36'b010011111100001100001000110111000011;
		finv_table[ 538] = 36'b010011111000110000011100110110111110;
		finv_table[ 539] = 36'b010011110101010100101010110110111010;
		finv_table[ 540] = 36'b010011110001111000110000110110110101;
		finv_table[ 541] = 36'b010011101110011100101000110110110001;
		finv_table[ 542] = 36'b010011101011000000011100110110101100;
		finv_table[ 543] = 36'b010011100111100100000100110110101000;
		finv_table[ 544] = 36'b010011100100000111100110110110100011;
		finv_table[ 545] = 36'b010011100000101010111100110110011111;
		finv_table[ 546] = 36'b010011011101100110101100110110011011;
		finv_table[ 547] = 36'b010011011001110001001110110110010110;
		finv_table[ 548] = 36'b010011010110101100101110110110010010;
		finv_table[ 549] = 36'b010011010011001111100000110110001101;
		finv_table[ 550] = 36'b010011001111110010001100110110001001;
		finv_table[ 551] = 36'b010011001100010100101100110110000100;
		finv_table[ 552] = 36'b010011001000110111000100110110000000;
		finv_table[ 553] = 36'b010011000101110001111100110101111100;
		finv_table[ 554] = 36'b010011000010010100000010110101110111;
		finv_table[ 555] = 36'b010010111110110110000000110101110011;
		finv_table[ 556] = 36'b010010111011110000100000110101101111;
		finv_table[ 557] = 36'b010010110111111001011100110101101010;
		finv_table[ 558] = 36'b010010110101001100011010110101100110;
		finv_table[ 559] = 36'b010010110001010101000100110101100001;
		finv_table[ 560] = 36'b010010101110001111000110110101011101;
		finv_table[ 561] = 36'b010010101010110000001100110101011001;
		finv_table[ 562] = 36'b010010100111101001111100110101010101;
		finv_table[ 563] = 36'b010010100100001010110010110101010000;
		finv_table[ 564] = 36'b010010100000101011011100110101001100;
		finv_table[ 565] = 36'b010010011101100100110100110101001000;
		finv_table[ 566] = 36'b010010011010000101010000110101000011;
		finv_table[ 567] = 36'b010010010110111110010110110100111111;
		finv_table[ 568] = 36'b010010010011011110100000110100111011;
		finv_table[ 569] = 36'b010010010000010111011000110100110111;
		finv_table[ 570] = 36'b010010001100110111001100110100110010;
		finv_table[ 571] = 36'b010010001001101111110100110100101110;
		finv_table[ 572] = 36'b010010000110001111011000110100101010;
		finv_table[ 573] = 36'b010010000011000111110000110100100110;
		finv_table[ 574] = 36'b010010000000000000000000110100100010;
		finv_table[ 575] = 36'b010001111100011111001010110100011101;
		finv_table[ 576] = 36'b010001111000111110001000110100011001;
		finv_table[ 577] = 36'b010001110110001111000010110100010101;
		finv_table[ 578] = 36'b010001110010101101110000110100010001;
		finv_table[ 579] = 36'b010001101111001100010110110100001100;
		finv_table[ 580] = 36'b010001101100011100111000110100001001;
		finv_table[ 581] = 36'b010001101000111011001110110100000100;
		finv_table[ 582] = 36'b010001100101011001010110110100000000;
		finv_table[ 583] = 36'b010001100010101001100110110011111100;
		finv_table[ 584] = 36'b010001011111000111011110110011111000;
		finv_table[ 585] = 36'b010001011011111110010110110011110100;
		finv_table[ 586] = 36'b010001011000011011111100110011101111;
		finv_table[ 587] = 36'b010001010101101011101110110011101100;
		finv_table[ 588] = 36'b010001010010001001000100110011100111;
		finv_table[ 589] = 36'b010001001110111111011010110011100011;
		finv_table[ 590] = 36'b010001001011110101101100110011011111;
		finv_table[ 591] = 36'b010001001000101011110010110011011011;
		finv_table[ 592] = 36'b010001000101001000100100110011010111;
		finv_table[ 593] = 36'b010001000010010111101100110011010011;
		finv_table[ 594] = 36'b010000111110110100001000110011001111;
		finv_table[ 595] = 36'b010000111011101001110000110011001011;
		finv_table[ 596] = 36'b010000111000111000100110110011000111;
		finv_table[ 597] = 36'b010000110101010100101000110011000011;
		finv_table[ 598] = 36'b010000110010001001111000110010111111;
		finv_table[ 599] = 36'b010000101110111111000000110010111011;
		finv_table[ 600] = 36'b010000101011110100000000110010110111;
		finv_table[ 601] = 36'b010000101000101000111000110010110011;
		finv_table[ 602] = 36'b010000100101011101101000110010101111;
		finv_table[ 603] = 36'b010000100010010010010000110010101011;
		finv_table[ 604] = 36'b010000011111000110110000110010100111;
		finv_table[ 605] = 36'b010000011011111011001000110010100011;
		finv_table[ 606] = 36'b010000011000101111011000110010011111;
		finv_table[ 607] = 36'b010000010101100011100000110010011011;
		finv_table[ 608] = 36'b010000010010110001000000110010010111;
		finv_table[ 609] = 36'b010000001111001011011000110010010011;
		finv_table[ 610] = 36'b010000001100011000101010110010001111;
		finv_table[ 611] = 36'b010000001000110010110000110010001011;
		finv_table[ 612] = 36'b010000000101111111110100110010000111;
		finv_table[ 613] = 36'b010000000010110011001010110010000011;
		finv_table[ 614] = 36'b010000000000000000000000110010000000;
		finv_table[ 615] = 36'b001111111100011001100010110001111011;
		finv_table[ 616] = 36'b001111111001100110001010110001111000;
		finv_table[ 617] = 36'b001111110101111111011000110001110011;
		finv_table[ 618] = 36'b001111110011100101011100110001110000;
		finv_table[ 619] = 36'b001111101111111110011010110001101100;
		finv_table[ 620] = 36'b001111101101001010100110110001101000;
		finv_table[ 621] = 36'b001111101001100011010000110001100100;
		finv_table[ 622] = 36'b001111100111001000111100110001100001;
		finv_table[ 623] = 36'b001111100011100001010110110001011100;
		finv_table[ 624] = 36'b001111100000101101000100110001011001;
		finv_table[ 625] = 36'b001111011101011110111100110001010101;
		finv_table[ 626] = 36'b001111011010101010100000110001010001;
		finv_table[ 627] = 36'b001111010111000010010100110001001101;
		finv_table[ 628] = 36'b001111010100100111011100110001001010;
		finv_table[ 629] = 36'b001111010000111111000000110001000101;
		finv_table[ 630] = 36'b001111001110001010000110110001000010;
		finv_table[ 631] = 36'b001111001011010101000100110000111110;
		finv_table[ 632] = 36'b001111001000000110000100110000111010;
		finv_table[ 633] = 36'b001111000100110110111110110000110110;
		finv_table[ 634] = 36'b001111000010000001101000110000110011;
		finv_table[ 635] = 36'b001110111110110010010000110000101111;
		finv_table[ 636] = 36'b001110111011111100101100110000101011;
		finv_table[ 637] = 36'b001110111000101101000010110000100111;
		finv_table[ 638] = 36'b001110110101110111010000110000100100;
		finv_table[ 639] = 36'b001110110010100111011000110000100000;
		finv_table[ 640] = 36'b001110101111110001011000110000011100;
		finv_table[ 641] = 36'b001110101100111011010000110000011001;
		finv_table[ 642] = 36'b001110101001101011000000110000010101;
		finv_table[ 643] = 36'b001110100110011010101000110000010001;
		finv_table[ 644] = 36'b001110100011100100001110110000001101;
		finv_table[ 645] = 36'b001110100000101101101010110000001010;
		finv_table[ 646] = 36'b001110011101110111000000110000000110;
		finv_table[ 647] = 36'b001110011010100110001010110000000010;
		finv_table[ 648] = 36'b001110010111010101001000101111111110;
		finv_table[ 649] = 36'b001110010100111000010010101111111011;
		finv_table[ 650] = 36'b001110010001100111000100101111110111;
		finv_table[ 651] = 36'b001110001110010101101010101111110011;
		finv_table[ 652] = 36'b001110001011111000100010101111110000;
		finv_table[ 653] = 36'b001110001000100110111100101111101100;
		finv_table[ 654] = 36'b001110000101101111011000101111101001;
		finv_table[ 655] = 36'b001110000010011101100000101111100101;
		finv_table[ 656] = 36'b001110000000000000000000101111100010;
		finv_table[ 657] = 36'b001101111100101101111000101111011110;
		finv_table[ 658] = 36'b001101111001110101111010101111011010;
		finv_table[ 659] = 36'b001101110110100011100100101111010110;
		finv_table[ 660] = 36'b001101110100000101101100101111010011;
		finv_table[ 661] = 36'b001101110000110011000010101111001111;
		finv_table[ 662] = 36'b001101101101111010101000101111001100;
		finv_table[ 663] = 36'b001101101011000010001000101111001000;
		finv_table[ 664] = 36'b001101101000001001100000101111000101;
		finv_table[ 665] = 36'b001101100101010000110000101111000001;
		finv_table[ 666] = 36'b001101100010010111111010101110111110;
		finv_table[ 667] = 36'b001101011111000100100010101110111010;
		finv_table[ 668] = 36'b001101011100001011011110101110110110;
		finv_table[ 669] = 36'b001101011001101100110000101110110011;
		finv_table[ 670] = 36'b001101010110011001000010101110101111;
		finv_table[ 671] = 36'b001101010011011111101000101110101100;
		finv_table[ 672] = 36'b001101010000100110001000101110101000;
		finv_table[ 673] = 36'b001101001101101100100000101110100101;
		finv_table[ 674] = 36'b001101001011001101010100101110100010;
		finv_table[ 675] = 36'b001101000111111000111100101110011110;
		finv_table[ 676] = 36'b001101000100111111000000101110011010;
		finv_table[ 677] = 36'b001101000010000100111100101110010111;
		finv_table[ 678] = 36'b001100111111001010110100101110010011;
		finv_table[ 679] = 36'b001100111100010000100010101110010000;
		finv_table[ 680] = 36'b001100111001010110001010101110001100;
		finv_table[ 681] = 36'b001100110110110110010100101110001001;
		finv_table[ 682] = 36'b001100110011100001000110101110000101;
		finv_table[ 683] = 36'b001100110001000001000100101110000010;
		finv_table[ 684] = 36'b001100101101101011100010101101111110;
		finv_table[ 685] = 36'b001100101011001011010100101101111011;
		finv_table[ 686] = 36'b001100101000010000010010101101111000;
		finv_table[ 687] = 36'b001100100101010101001010101101110100;
		finv_table[ 688] = 36'b001100100010011001111000101101110001;
		finv_table[ 689] = 36'b001100011111011110100010101101101101;
		finv_table[ 690] = 36'b001100011100111101110110101101101010;
		finv_table[ 691] = 36'b001100011001100111100000101101100110;
		finv_table[ 692] = 36'b001100010111000110101000101101100011;
		finv_table[ 693] = 36'b001100010100001010110100101101100000;
		finv_table[ 694] = 36'b001100010001001110111000101101011100;
		finv_table[ 695] = 36'b001100001110101101110000101101011001;
		finv_table[ 696] = 36'b001100001011110001101000101101010110;
		finv_table[ 697] = 36'b001100001000110101011010101101010010;
		finv_table[ 698] = 36'b001100000101111001000100101101001111;
		finv_table[ 699] = 36'b001100000011010111100000101101001100;
		finv_table[ 700] = 36'b001100000000011010111100101101001000;
		finv_table[ 701] = 36'b001011111101011110010010101101000101;
		finv_table[ 702] = 36'b001011111010100001100000101101000001;
		finv_table[ 703] = 36'b001011110111111111100110101100111110;
		finv_table[ 704] = 36'b001011110101000010100100101100111011;
		finv_table[ 705] = 36'b001011110010100000100000101100111000;
		finv_table[ 706] = 36'b001011101111100011010010101100110100;
		finv_table[ 707] = 36'b001011101100100101111100101100110001;
		finv_table[ 708] = 36'b001011101010000011100100101100101110;
		finv_table[ 709] = 36'b001011100111000110000010101100101010;
		finv_table[ 710] = 36'b001011100100001000011000101100100111;
		finv_table[ 711] = 36'b001011100001100101101110101100100100;
		finv_table[ 712] = 36'b001011011110100111110110101100100000;
		finv_table[ 713] = 36'b001011011100000101000000101100011101;
		finv_table[ 714] = 36'b001011011001000110111010101100011010;
		finv_table[ 715] = 36'b001011010110100011111000101100010111;
		finv_table[ 716] = 36'b001011010011100101100100101100010011;
		finv_table[ 717] = 36'b001011010001000010010110101100010000;
		finv_table[ 718] = 36'b001011001110000011110100101100001101;
		finv_table[ 719] = 36'b001011001011100000011010101100001010;
		finv_table[ 720] = 36'b001011001000100001101010101100000110;
		finv_table[ 721] = 36'b001011000101100010110100101100000011;
		finv_table[ 722] = 36'b001011000011011010011000101100000000;
		finv_table[ 723] = 36'b001011000000011011010100101011111101;
		finv_table[ 724] = 36'b001010111101011100001000101011111001;
		finv_table[ 725] = 36'b001010111010111000001010101011110110;
		finv_table[ 726] = 36'b001010110111111000110000101011110011;
		finv_table[ 727] = 36'b001010110101101111111110101011110000;
		finv_table[ 728] = 36'b001010110010010100111100101011101100;
		finv_table[ 729] = 36'b001010110000001100000000101011101010;
		finv_table[ 730] = 36'b001010101101001100001010101011100110;
		finv_table[ 731] = 36'b001010101010001100001100101011100011;
		finv_table[ 732] = 36'b001010101000000011000000101011100000;
		finv_table[ 733] = 36'b001010100101000010110110101011011101;
		finv_table[ 734] = 36'b001010100010000010100100101011011001;
		finv_table[ 735] = 36'b001010011111111001001000101011010111;
		finv_table[ 736] = 36'b001010011100111000101010101011010011;
		finv_table[ 737] = 36'b001010011001111000000010101011010000;
		finv_table[ 738] = 36'b001010010111101110011000101011001101;
		finv_table[ 739] = 36'b001010010100101101100010101011001010;
		finv_table[ 740] = 36'b001010010010001000001100101011000111;
		finv_table[ 741] = 36'b001010001111100010101100101011000100;
		finv_table[ 742] = 36'b001010001100100001100010101011000000;
		finv_table[ 743] = 36'b001010001001111011111000101010111101;
		finv_table[ 744] = 36'b001010000111010110001000101010111010;
		finv_table[ 745] = 36'b001010000100110000010010101010110111;
		finv_table[ 746] = 36'b001010000010001010010110101010110100;
		finv_table[ 747] = 36'b001001111111001000101000101010110001;
		finv_table[ 748] = 36'b001001111100100010100010101010101110;
		finv_table[ 749] = 36'b001001111010011000000000101010101011;
		finv_table[ 750] = 36'b001001110110111010010010101010100111;
		finv_table[ 751] = 36'b001001110100101111100100101010100101;
		finv_table[ 752] = 36'b001001110010001001000110101010100010;
		finv_table[ 753] = 36'b001001101111000110110000101010011110;
		finv_table[ 754] = 36'b001001101100111011110100101010011100;
		finv_table[ 755] = 36'b001001101001111001010000101010011000;
		finv_table[ 756] = 36'b001001100111010010011000101010010101;
		finv_table[ 757] = 36'b001001100100101011011010101010010010;
		finv_table[ 758] = 36'b001001100010000100010110101010001111;
		finv_table[ 759] = 36'b001001011111011101001100101010001100;
		finv_table[ 760] = 36'b001001011100110101111100101010001001;
		finv_table[ 761] = 36'b001001011010001110100110101010000110;
		finv_table[ 762] = 36'b001001010111100111001010101010000011;
		finv_table[ 763] = 36'b001001010100111111101000101010000000;
		finv_table[ 764] = 36'b001001010010011000000000101001111101;
		finv_table[ 765] = 36'b001001001111110000010010101001111010;
		finv_table[ 766] = 36'b001001001101001000011110101001110111;
		finv_table[ 767] = 36'b001001001010000100100100101001110100;
		finv_table[ 768] = 36'b001001000111111000100100101001110001;
		finv_table[ 769] = 36'b001001000101010000100000101001101110;
		finv_table[ 770] = 36'b001001000010101000010100101001101011;
		finv_table[ 771] = 36'b001001000000000000000010101001101000;
		finv_table[ 772] = 36'b001000111101010111101000101001100101;
		finv_table[ 773] = 36'b001000111011001011010000101001100011;
		finv_table[ 774] = 36'b001000111000000110100110101001011111;
		finv_table[ 775] = 36'b001000110101011101111100101001011100;
		finv_table[ 776] = 36'b001000110011010001010100101001011010;
		finv_table[ 777] = 36'b001000110000001100010110101001010110;
		finv_table[ 778] = 36'b001000101101111111100010101001010100;
		finv_table[ 779] = 36'b001000101011010110100000101001010001;
		finv_table[ 780] = 36'b001000101000101101011000101001001110;
		finv_table[ 781] = 36'b001000100110000100001100101001001011;
		finv_table[ 782] = 36'b001000100011011010110110101001001000;
		finv_table[ 783] = 36'b001000100001001101101100101001000101;
		finv_table[ 784] = 36'b001000011110100100001100101001000010;
		finv_table[ 785] = 36'b001000011011111010100110101000111111;
		finv_table[ 786] = 36'b001000011001010000111010101000111100;
		finv_table[ 787] = 36'b001000010110100111001000101000111001;
		finv_table[ 788] = 36'b001000010100011001100100101000110111;
		finv_table[ 789] = 36'b001000010001010011010000101000110011;
		finv_table[ 790] = 36'b001000001111000101100100101000110001;
		finv_table[ 791] = 36'b001000001100110111110000101000101110;
		finv_table[ 792] = 36'b001000001001110001001000101000101011;
		finv_table[ 793] = 36'b001000000111100011001100101000101000;
		finv_table[ 794] = 36'b001000000100111000110000101000100101;
		finv_table[ 795] = 36'b001000000010001110001110101000100010;
		finv_table[ 796] = 36'b001000000000000000000000101000100000;
		finv_table[ 797] = 36'b000111111101010101010100101000011101;
		finv_table[ 798] = 36'b000111111010101010011110101000011010;
		finv_table[ 799] = 36'b000111111000011100000100101000010111;
		finv_table[ 800] = 36'b000111110101110001000100101000010100;
		finv_table[ 801] = 36'b000111110011000101111110101000010001;
		finv_table[ 802] = 36'b000111110000110111010100101000001111;
		finv_table[ 803] = 36'b000111101110001100000010101000001100;
		finv_table[ 804] = 36'b000111101011111101001110101000001001;
		finv_table[ 805] = 36'b000111101000110101001010101000000110;
		finv_table[ 806] = 36'b000111100111000010110010101000000100;
		finv_table[ 807] = 36'b000111100011111010100010101000000000;
		finv_table[ 808] = 36'b000111100001101011011010100111111110;
		finv_table[ 809] = 36'b000111011111011100001100100111111011;
		finv_table[ 810] = 36'b000111011100010011100110100111111000;
		finv_table[ 811] = 36'b000111011010100000111010100111110110;
		finv_table[ 812] = 36'b000111010111110100110100100111110011;
		finv_table[ 813] = 36'b000111010101001000100100100111110000;
		finv_table[ 814] = 36'b000111010010011100010000100111101101;
		finv_table[ 815] = 36'b000111010000101001010100100111101011;
		finv_table[ 816] = 36'b000111001101100000000110100111100111;
		finv_table[ 817] = 36'b000111001011010000010000100111100101;
		finv_table[ 818] = 36'b000111001001000000010110100111100010;
		finv_table[ 819] = 36'b000111000110010011100100100111011111;
		finv_table[ 820] = 36'b000111000100000011100000100111011101;
		finv_table[ 821] = 36'b000111000001010110100010100111011010;
		finv_table[ 822] = 36'b000110111111000110010100100111010111;
		finv_table[ 823] = 36'b000110111100011001001010100111010100;
		finv_table[ 824] = 36'b000110111010001000110010100111010010;
		finv_table[ 825] = 36'b000110110111011011011100100111001111;
		finv_table[ 826] = 36'b000110110101001010111010100111001100;
		finv_table[ 827] = 36'b000110110010111010010010100111001010;
		finv_table[ 828] = 36'b000110110000001100101100100111000111;
		finv_table[ 829] = 36'b000110101101111011111010100111000100;
		finv_table[ 830] = 36'b000110101011001110000110100111000001;
		finv_table[ 831] = 36'b000110101000111101001100100110111111;
		finv_table[ 832] = 36'b000110100110101100001010100110111100;
		finv_table[ 833] = 36'b000110100011111110000100100110111001;
		finv_table[ 834] = 36'b000110100001101100111100100110110111;
		finv_table[ 835] = 36'b000110011110111110101000100110110100;
		finv_table[ 836] = 36'b000110011100101101010110100110110001;
		finv_table[ 837] = 36'b000110011010011011111100100110101111;
		finv_table[ 838] = 36'b000110011000001010011110100110101100;
		finv_table[ 839] = 36'b000110010101011011110100100110101001;
		finv_table[ 840] = 36'b000110010011001010001100100110100111;
		finv_table[ 841] = 36'b000110010000111000100000100110100100;
		finv_table[ 842] = 36'b000110001110001001100100100110100001;
		finv_table[ 843] = 36'b000110001011110111101100100110011111;
		finv_table[ 844] = 36'b000110001001100101110000100110011100;
		finv_table[ 845] = 36'b000110000110110110100010100110011001;
		finv_table[ 846] = 36'b000110000100100100011100100110010111;
		finv_table[ 847] = 36'b000110000010010010010000100110010100;
		finv_table[ 848] = 36'b000110000000000000000000100110010010;
		finv_table[ 849] = 36'b000101111101101101101100100110001111;
		finv_table[ 850] = 36'b000101111010111110000000100110001100;
		finv_table[ 851] = 36'b000101111000101011100000100110001010;
		finv_table[ 852] = 36'b000101110110011000111110100110000111;
		finv_table[ 853] = 36'b000101110100000110010100100110000101;
		finv_table[ 854] = 36'b000101110001010110010000100110000010;
		finv_table[ 855] = 36'b000101101111100000110100100110000000;
		finv_table[ 856] = 36'b000101101100110000100100100101111101;
		finv_table[ 857] = 36'b000101101010011101101000100101111010;
		finv_table[ 858] = 36'b000101101000001010100100100101111000;
		finv_table[ 859] = 36'b000101100101011010000100100101110101;
		finv_table[ 860] = 36'b000101100011100100010100100101110011;
		finv_table[ 861] = 36'b000101100000110011100100100101110000;
		finv_table[ 862] = 36'b000101011110111101101100100101101110;
		finv_table[ 863] = 36'b000101011100001100110100100101101011;
		finv_table[ 864] = 36'b000101011001111001010010100101101000;
		finv_table[ 865] = 36'b000101010111100101101110100101100110;
		finv_table[ 866] = 36'b000101010101010010000100100101100011;
		finv_table[ 867] = 36'b000101010010111110010100100101100001;
		finv_table[ 868] = 36'b000101010000101010100000100101011110;
		finv_table[ 869] = 36'b000101001101111001000010100101011011;
		finv_table[ 870] = 36'b000101001100000010101100100101011001;
		finv_table[ 871] = 36'b000101001001101110101000100101010111;
		finv_table[ 872] = 36'b000101000110111100111000100101010100;
		finv_table[ 873] = 36'b000101000101000110010100100101010010;
		finv_table[ 874] = 36'b000101000010010100011000100101001111;
		finv_table[ 875] = 36'b000101000000011101101100100101001101;
		finv_table[ 876] = 36'b000100111101101011100100100101001010;
		finv_table[ 877] = 36'b000100111011110100110000100101001000;
		finv_table[ 878] = 36'b000100111001000010011100100101000101;
		finv_table[ 879] = 36'b000100110110101101110010100101000010;
		finv_table[ 880] = 36'b000100110100110110110000100101000000;
		finv_table[ 881] = 36'b000100110010100001111100100100111110;
		finv_table[ 882] = 36'b000100101111101111010000100100111011;
		finv_table[ 883] = 36'b000100101101111000000100100100111001;
		finv_table[ 884] = 36'b000100101011000101001100100100110110;
		finv_table[ 885] = 36'b000100101001001101111000100100110100;
		finv_table[ 886] = 36'b000100100110111000101010100100110001;
		finv_table[ 887] = 36'b000100100100100011011000100100101111;
		finv_table[ 888] = 36'b000100100010001101111110100100101100;
		finv_table[ 889] = 36'b000100011111111000100010100100101010;
		finv_table[ 890] = 36'b000100011101100011000000100100100111;
		finv_table[ 891] = 36'b000100011011001101011000100100100101;
		finv_table[ 892] = 36'b000100011001010101101000100100100011;
		finv_table[ 893] = 36'b000100010110100001111100100100100000;
		finv_table[ 894] = 36'b000100010100101010000100100100011110;
		finv_table[ 895] = 36'b000100010001110110001000100100011011;
		finv_table[ 896] = 36'b000100001111111110001000100100011001;
		finv_table[ 897] = 36'b000100001101101000000100100100010110;
		finv_table[ 898] = 36'b000100001011101111111100100100010100;
		finv_table[ 899] = 36'b000100001000111011101010100100010001;
		finv_table[ 900] = 36'b000100000111000011011010100100001111;
		finv_table[ 901] = 36'b000100000100001110111100100100001100;
		finv_table[ 902] = 36'b000100000010010110100100100100001010;
		finv_table[ 903] = 36'b000100000000000000000000100100001000;
		finv_table[ 904] = 36'b000011111110000111100000100100000110;
		finv_table[ 905] = 36'b000011111011010010101100100100000011;
		finv_table[ 906] = 36'b000011111001011010000100100100000001;
		finv_table[ 907] = 36'b000011110111000011001100100011111110;
		finv_table[ 908] = 36'b000011110100101100010000100011111100;
		finv_table[ 909] = 36'b000011110010110011011100100011111010;
		finv_table[ 910] = 36'b000011110000011100010110100011110111;
		finv_table[ 911] = 36'b000011101110000101001100100011110101;
		finv_table[ 912] = 36'b000011101011101101111010100011110010;
		finv_table[ 913] = 36'b000011101001010110100110100011110000;
		finv_table[ 914] = 36'b000011100111011101011110100011101110;
		finv_table[ 915] = 36'b000011100101000101111110100011101011;
		finv_table[ 916] = 36'b000011100011001100110000100011101001;
		finv_table[ 917] = 36'b000011100000010110110010100011100110;
		finv_table[ 918] = 36'b000011011110011101011000100011100100;
		finv_table[ 919] = 36'b000011011100100011111110100011100010;
		finv_table[ 920] = 36'b000011011001101101101110100011011111;
		finv_table[ 921] = 36'b000011010111110100001000100011011101;
		finv_table[ 922] = 36'b000011010101111010100010100011011011;
		finv_table[ 923] = 36'b000011010011000100000000100011011000;
		finv_table[ 924] = 36'b000011010001001010001110100011010110;
		finv_table[ 925] = 36'b000011001111010000011100100011010100;
		finv_table[ 926] = 36'b000011001100011001101000100011010001;
		finv_table[ 927] = 36'b000011001010111110001010100011010000;
		finv_table[ 928] = 36'b000011001000000111001010100011001101;
		finv_table[ 929] = 36'b000011000110001101000100100011001011;
		finv_table[ 930] = 36'b000011000011110100011100100011001000;
		finv_table[ 931] = 36'b000011000001111010010000100011000110;
		finv_table[ 932] = 36'b000010111111100001011100100011000100;
		finv_table[ 933] = 36'b000010111101001000100010100011000001;
		finv_table[ 934] = 36'b000010111011001110001100100010111111;
		finv_table[ 935] = 36'b000010111001010011101110100010111101;
		finv_table[ 936] = 36'b000010110110011011111110100010111010;
		finv_table[ 937] = 36'b000010110101000000000100100010111001;
		finv_table[ 938] = 36'b000010110010001000001000100010110110;
		finv_table[ 939] = 36'b000010110000001101011100100010110100;
		finv_table[ 940] = 36'b000010101110010010101100100010110010;
		finv_table[ 941] = 36'b000010101011111001001010100010101111;
		finv_table[ 942] = 36'b000010101001111110010100100010101101;
		finv_table[ 943] = 36'b000010100111100100101000100010101011;
		finv_table[ 944] = 36'b000010100101001010111000100010101000;
		finv_table[ 945] = 36'b000010100011001111110100100010100110;
		finv_table[ 946] = 36'b000010100001010100101100100010100100;
		finv_table[ 947] = 36'b000010011110111010101100100010100010;
		finv_table[ 948] = 36'b000010011100100000101010100010011111;
		finv_table[ 949] = 36'b000010011010100101010100100010011101;
		finv_table[ 950] = 36'b000010011000101001111110100010011011;
		finv_table[ 951] = 36'b000010010110001111101000100010011001;
		finv_table[ 952] = 36'b000010010100010100001000100010010111;
		finv_table[ 953] = 36'b000010010001111001101110100010010100;
		finv_table[ 954] = 36'b000010001111111110000100100010010010;
		finv_table[ 955] = 36'b000010001101100011011110100010010000;
		finv_table[ 956] = 36'b000010001011100111101110100010001110;
		finv_table[ 957] = 36'b000010001001101011111010100010001100;
		finv_table[ 958] = 36'b000010000111010001000100100010001001;
		finv_table[ 959] = 36'b000010000101010101001000100010000111;
		finv_table[ 960] = 36'b000010000010111010001000100010000101;
		finv_table[ 961] = 36'b000010000000111110000100100010000011;
		finv_table[ 962] = 36'b000001111111000001111100100010000001;
		finv_table[ 963] = 36'b000001111100100110101110100001111110;
		finv_table[ 964] = 36'b000001111010001011011000100001111100;
		finv_table[ 965] = 36'b000001111000101110001010100001111010;
		finv_table[ 966] = 36'b000001110110010010101100100001111000;
		finv_table[ 967] = 36'b000001110100010110010000100001110110;
		finv_table[ 968] = 36'b000001110001111010101000100001110011;
		finv_table[ 969] = 36'b000001101111111110000100100001110001;
		finv_table[ 970] = 36'b000001101110000001011100100001101111;
		finv_table[ 971] = 36'b000001101011100101100100100001101101;
		finv_table[ 972] = 36'b000001101001101000110100100001101011;
		finv_table[ 973] = 36'b000001100111101100000000100001101001;
		finv_table[ 974] = 36'b000001100101001111111010100001100110;
		finv_table[ 975] = 36'b000001100011010011000000100001100100;
		finv_table[ 976] = 36'b000001100001010101111110100001100010;
		finv_table[ 977] = 36'b000001011111011000111100100001100000;
		finv_table[ 978] = 36'b000001011100111100100000100001011110;
		finv_table[ 979] = 36'b000001011010111111010100100001011100;
		finv_table[ 980] = 36'b000001011001000010000100100001011010;
		finv_table[ 981] = 36'b000001010110100101011100100001010111;
		finv_table[ 982] = 36'b000001010100101000000100100001010101;
		finv_table[ 983] = 36'b000001010010101010101000100001010011;
		finv_table[ 984] = 36'b000001010000101101001000100001010001;
		finv_table[ 985] = 36'b000001001110010000001100100001001111;
		finv_table[ 986] = 36'b000001001100110001111110100001001101;
		finv_table[ 987] = 36'b000001001010010100110110100001001011;
		finv_table[ 988] = 36'b000001000111110111101010100001001000;
		finv_table[ 989] = 36'b000001000110011001010100100001000111;
		finv_table[ 990] = 36'b000001000011111011111100100001000100;
		finv_table[ 991] = 36'b000001000001111110000010100001000010;
		finv_table[ 992] = 36'b000001000000000000000000100001000000;
		finv_table[ 993] = 36'b000000111110000001111110100000111110;
		finv_table[ 994] = 36'b000000111100000011110100100000111100;
		finv_table[ 995] = 36'b000000111001100110000110100000111010;
		finv_table[ 996] = 36'b000000111000000111011010100000111000;
		finv_table[ 997] = 36'b000000110101101001100000100000110110;
		finv_table[ 998] = 36'b000000110011101011001000100000110100;
		finv_table[ 999] = 36'b000000110001001101000110100000110001;
		finv_table[1000] = 36'b000000101111101110001110100000110000;
		finv_table[1001] = 36'b000000101101010000000000100000101101;
		finv_table[1002] = 36'b000000101011110001000010100000101100;
		finv_table[1003] = 36'b000000101001010010101100100000101001;
		finv_table[1004] = 36'b000000100111010011111100100000100111;
		finv_table[1005] = 36'b000000100101010101001000100000100101;
		finv_table[1006] = 36'b000000100011010110010000100000100011;
		finv_table[1007] = 36'b000000100001010111010100100000100001;
		finv_table[1008] = 36'b000000011111011000010100100000011111;
		finv_table[1009] = 36'b000000011100111001100000100000011101;
		finv_table[1010] = 36'b000000011011011010001010100000011011;
		finv_table[1011] = 36'b000000011000111011001000100000011001;
		finv_table[1012] = 36'b000000010111011011101110100000010111;
		finv_table[1013] = 36'b000000010100111100100100100000010101;
		finv_table[1014] = 36'b000000010010111101001100100000010011;
		finv_table[1015] = 36'b000000010000111101110000100000010001;
		finv_table[1016] = 36'b000000001111011110001010100000001111;
		finv_table[1017] = 36'b000000001100111110101100100000001101;
		finv_table[1018] = 36'b000000001010111111000100100000001011;
		finv_table[1019] = 36'b000000001000111111011000100000001001;
		finv_table[1020] = 36'b000000000110111111101000100000000111;
		finv_table[1021] = 36'b000000000100111111110100100000000101;
		finv_table[1022] = 36'b000000000010111111111100100000000011;
		finv_table[1023] = 36'b000000000001000000000000100000000001;
	end
endmodule

`default_nettype wire