`default_nettype wire
module sqrt (
	input logic [31:0]  x,
  output logic [31:0] y,
  //output logic        ovf,
  input logic       clk,
  input logic       rstn
);
	// step1
	wire [ 7:0] exp_x = x[30:23];
	wire [ 7:0] exp_x_unbiased = {exp_x - 8'd127};
	wire [ 7:0] exp_y_unbiased = {exp_x_unbiased[7],exp_x_unbiased[7:1]};// >> 1 ;
	wire [ 7:0] exp_y = exp_y_unbiased + 8'd127;
	wire [ 9:0] addr = {~x[23],x[22:14]};

	// step2
	wire [35:0] dout;
	sqrt_table sqrt_table1(addr_reg, dout, clk, rstn);

	wire [12:0] dx = (x_reg1[23]) ? {1'b0, 8'b0,1'b0,x_reg1[13:11]} : {1'b0, 7'b0,1'b0,x_reg1[14:11]} ;//(x[23]) ? : x[12:0];
	wire [12:0] gradient = dout[12:0];
	wire [26:0] dy_calc = gradient * dx;

	// step3
	wire [22:0] constant = dout_reg[35:13];
	wire [22:0] tmp =  constant + dy_calc_reg[26:4];// + dy_calc[26:4];
	wire [22:0] frac_y = {tmp[21:0],1'b0};

	assign y = (x_reg2[30:23] == 8'b0) ? 32'b0 : {1'b0 , exp_y_reg2, frac_y};

	// reg
	logic [31:0] x_reg1, x_reg2;
	logic [35:0] dout_reg;
	logic [ 7:0] exp_y_reg1, exp_y_reg2;
	logic [ 9:0] addr_reg;
	logic [26:0] dy_calc_reg;
	always_ff @( posedge clk ) begin
		if (~rstn) begin
			x_reg1 <= 32'b0;
			x_reg2 <= 32'b0;
			dout_reg <= 36'b0;
			exp_y_reg1 <= 8'b0;
			exp_y_reg2 <= 8'b0;
			addr_reg <= 10'b0;
			dy_calc_reg <= 27'b0;
		end else begin
			x_reg1 <= x;
			x_reg2 <= x_reg1;
			dout_reg <= dout;
			exp_y_reg1 <= exp_y;
			exp_y_reg2 <= exp_y_reg1;
			addr_reg <= addr;
			dy_calc_reg <= dy_calc;
		end
	end
endmodule

module sqrt_table (
	input		logic [ 9:0]	addr,
	output	logic  [35:0] dout,
	input 	logic 				clk,
	input 	logic 				rstn
);
	(*ram_style = "BLOCK"*) logic [35:0] sqrt_table [1023:0];
	always_comb begin
		dout = sqrt_table[addr];
	end
	initial begin
	 $readmemb("some_input.mem",sqrt_table);
		/*sqrt_table[   0] = 36'b10000000000110000000001_0111111111101;
		sqrt_table[   1] = 36'b100000000100100000100110111111110111;
		sqrt_table[   2] = 36'b100000000111100001101110111111110001;
		sqrt_table[   3] = 36'b100000001010011000101010111111101011;
		sqrt_table[   4] = 36'b100000001101011010111010111111100101;
		sqrt_table[   5] = 36'b100000010000011101101110111111011111;
		sqrt_table[   6] = 36'b100000010011100001000110111111011001;
		sqrt_table[   7] = 36'b100000010110001111010000111111010100;
		sqrt_table[   8] = 36'b100000011001011110101010111111001101;
		sqrt_table[   9] = 36'b100000011100001101110110111111001000;
		sqrt_table[  10] = 36'b100000011111010011011110111111000010;
		sqrt_table[  11] = 36'b100000100010001110101000111110111100;
		sqrt_table[  12] = 36'b100000100101001010010110111110110111;
		sqrt_table[  13] = 36'b100000101000000110100110111110110001;
		sqrt_table[  14] = 36'b100000101011000011010110111110101011;
		sqrt_table[  15] = 36'b100000101110000000101010111110100110;
		sqrt_table[  16] = 36'b100000110000110011010100111110100000;
		sqrt_table[  17] = 36'b100000110011111100111000111110011010;
		sqrt_table[  18] = 36'b100000110110110000100100111110010101;
		sqrt_table[  19] = 36'b100000111001100100101110111110010000;
		sqrt_table[  20] = 36'b100000111100100100101010111110001010;
		sqrt_table[  21] = 36'b100000111111100101001010111110000100;
		sqrt_table[  22] = 36'b100001000010011010110110111101111111;
		sqrt_table[  23] = 36'b100001000101010001000000111101111010;
		sqrt_table[  24] = 36'b100001001000010011000100111101110100;
		sqrt_table[  25] = 36'b100001001011001010010000111101101111;
		sqrt_table[  26] = 36'b100001001110000001111010111101101001;
		sqrt_table[  27] = 36'b100001010000111010000110111101100100;
		sqrt_table[  28] = 36'b100001010011110010110000111101011111;
		sqrt_table[  29] = 36'b100001010110100000010110111101011010;
		sqrt_table[  30] = 36'b100001011001100101100110111101010100;
		sqrt_table[  31] = 36'b100001011100011111110000111101001111;
		sqrt_table[  32] = 36'b100001011111001110110010111101001010;
		sqrt_table[  33] = 36'b100001100010001001111100111101000100;
		sqrt_table[  34] = 36'b100001100101000101101000111100111111;
		sqrt_table[  35] = 36'b100001100111110110000010111100111010;
		sqrt_table[  36] = 36'b100001101010100110111010111100110101;
		sqrt_table[  37] = 36'b100001101101100100000100111100110000;
		sqrt_table[  38] = 36'b100001110000100001101110111100101010;
		sqrt_table[  39] = 36'b100001110011001000001000111100100110;
		sqrt_table[  40] = 36'b100001110110000110110010111100100000;
		sqrt_table[  41] = 36'b100001111000111001111110111100011011;
		sqrt_table[  42] = 36'b100001111011111001101010111100010110;
		sqrt_table[  43] = 36'b100001111110100001110100111100010001;
		sqrt_table[  44] = 36'b100010000001010110011100111100001100;
		sqrt_table[  45] = 36'b100010000100010111101000111100000111;
		sqrt_table[  46] = 36'b100010000111000001000100111100000010;
		sqrt_table[  47] = 36'b100010001001110111000110111011111101;
		sqrt_table[  48] = 36'b100010001100100001011010111011111001;
		sqrt_table[  49] = 36'b100010001111100100100100111011110011;
		sqrt_table[  50] = 36'b100010010010001111110010111011101111;
		sqrt_table[  51] = 36'b100010010101000111101110111011101010;
		sqrt_table[  52] = 36'b100010010111110011110100111011100101;
		sqrt_table[  53] = 36'b100010011010101100101000111011100000;
		sqrt_table[  54] = 36'b100010011101011001100100111011011011;
		sqrt_table[  55] = 36'b100010100000010011011000111011010110;
		sqrt_table[  56] = 36'b100010100011000001001110111011010010;
		sqrt_table[  57] = 36'b100010100101101111100000111011001101;
		sqrt_table[  58] = 36'b100010101000101010101010111011001000;
		sqrt_table[  59] = 36'b100010101011001101010100111011000100;
		sqrt_table[  60] = 36'b100010101110001001011010111010111111;
		sqrt_table[  61] = 36'b100010110000111001011100111010111010;
		sqrt_table[  62] = 36'b100010110011101001111010111010110101;
		sqrt_table[  63] = 36'b100010110110001110001100111010110001;
		sqrt_table[  64] = 36'b100010111001001100001010111010101100;
		sqrt_table[  65] = 36'b100010111011111101111010111010100111;
		sqrt_table[  66] = 36'b100010111110100011011100111010100011;
		sqrt_table[  67] = 36'b100011000001010110000100111010011110;
		sqrt_table[  68] = 36'b100011000100001001001010111010011010;
		sqrt_table[  69] = 36'b100011000110101111110100111010010101;
		sqrt_table[  70] = 36'b100011001001110000101010111010010000;
		sqrt_table[  71] = 36'b100011001100001011010010111010001100;
		sqrt_table[  72] = 36'b100011001111000000001000111010001000;
		sqrt_table[  73] = 36'b100011010001110101011010111010000011;
		sqrt_table[  74] = 36'b100011010100011110000110111001111111;
		sqrt_table[  75] = 36'b100011010111000111001110111001111010;
		sqrt_table[  76] = 36'b100011011001111101110110111001110110;
		sqrt_table[  77] = 36'b100011011100100111110000111001110001;
		sqrt_table[  78] = 36'b100011011111010010001010111001101101;
		sqrt_table[  79] = 36'b100011100010001010000010111001101000;
		sqrt_table[  80] = 36'b100011100100101000000010111001100100;
		sqrt_table[  81] = 36'b100011100111100000110100111001100000;
		sqrt_table[  82] = 36'b100011101001111111100100111001011100;
		sqrt_table[  83] = 36'b100011101100111001001110111001010111;
		sqrt_table[  84] = 36'b100011101111011000101100111001010011;
		sqrt_table[  85] = 36'b100011110010010011001110111001001110;
		sqrt_table[  86] = 36'b100011110100110011011110111001001010;
		sqrt_table[  87] = 36'b100011110111100001011110111001000110;
		sqrt_table[  88] = 36'b100011111010001111111010111001000010;
		sqrt_table[  89] = 36'b100011111100111110101100111000111101;
		sqrt_table[  90] = 36'b100011111111100000011100111000111001;
		sqrt_table[  91] = 36'b100100000010010000001000111000110101;
		sqrt_table[  92] = 36'b100100000100110010101000111000110001;
		sqrt_table[  93] = 36'b100100000111100011000010111000101101;
		sqrt_table[  94] = 36'b100100001010010011111010111000101000;
		sqrt_table[  95] = 36'b100100001100101001111000111000100101;
		sqrt_table[  96] = 36'b100100001111101001001110111000100000;
		sqrt_table[  97] = 36'b100100010010001101100110111000011100;
		sqrt_table[  98] = 36'b100100010100110010011000111000011000;
		sqrt_table[  99] = 36'b100100010111010111011110111000010100;
		sqrt_table[ 100] = 36'b100100011001111100111110111000010000;
		sqrt_table[ 101] = 36'b100100011100110000101100111000001100;
		sqrt_table[ 102] = 36'b100100011111010110111100111000001000;
		sqrt_table[ 103] = 36'b100100100001111101100100111000000100;
		sqrt_table[ 104] = 36'b100100100100100100100100111000000000;
		sqrt_table[ 105] = 36'b100100100111001011111100110111111100;
		sqrt_table[ 106] = 36'b100100101010000001101000110111110111;
		sqrt_table[ 107] = 36'b100100101100011011110010110111110100;
		sqrt_table[ 108] = 36'b100100101111000100010010110111110000;
		sqrt_table[ 109] = 36'b100100110001101101001010110111101100;
		sqrt_table[ 110] = 36'b100100110100001000010010110111101000;
		sqrt_table[ 111] = 36'b100100110111000000000100110111100100;
		sqrt_table[ 112] = 36'b100100111001011011111000110111100000;
		sqrt_table[ 113] = 36'b100100111100000110010000110111011100;
		sqrt_table[ 114] = 36'b100100111110110001000000110111011000;
		sqrt_table[ 115] = 36'b100101000001001101111000110111010100;
		sqrt_table[ 116] = 36'b100101000011111001011000110111010000;
		sqrt_table[ 117] = 36'b100101000110100101010000110111001100;
		sqrt_table[ 118] = 36'b100101001001000011001000110111001001;
		sqrt_table[ 119] = 36'b100101001011100001011010110111000101;
		sqrt_table[ 120] = 36'b100101001110001110011010110111000001;
		sqrt_table[ 121] = 36'b100101010000111011110010110110111101;
		sqrt_table[ 122] = 36'b100101010011011011000000110110111001;
		sqrt_table[ 123] = 36'b100101010101111010101010110110110110;
		sqrt_table[ 124] = 36'b100101011000011010100110110110110010;
		sqrt_table[ 125] = 36'b100101011011001001011110110110101110;
		sqrt_table[ 126] = 36'b100101011101101010000110110110101010;
		sqrt_table[ 127] = 36'b100101100000001011000110110110100111;
		sqrt_table[ 128] = 36'b100101100010111011000110110110100011;
		sqrt_table[ 129] = 36'b100101100101001110000100110110011111;
		sqrt_table[ 130] = 36'b100101100111111110110100110110011011;
		sqrt_table[ 131] = 36'b100101101010010010011100110110011000;
		sqrt_table[ 132] = 36'b100101101101000011111100110110010100;
		sqrt_table[ 133] = 36'b100101101111011000001010110110010001;
		sqrt_table[ 134] = 36'b100101110010001010011010110110001101;
		sqrt_table[ 135] = 36'b100101110100101110001100110110001001;
		sqrt_table[ 136] = 36'b100101110111000011010110110110000110;
		sqrt_table[ 137] = 36'b100101111001100111110000110110000010;
		sqrt_table[ 138] = 36'b100101111100001100100010110101111110;
		sqrt_table[ 139] = 36'b100101111110110001101000110101111011;
		sqrt_table[ 140] = 36'b100110000001010111001000110101110111;
		sqrt_table[ 141] = 36'b100110000011101101110110110101110100;
		sqrt_table[ 142] = 36'b100110000110010011111110110101110000;
		sqrt_table[ 143] = 36'b100110001000101011010100110101101101;
		sqrt_table[ 144] = 36'b100110001011100001010100110101101001;
		sqrt_table[ 145] = 36'b100110001101111001010010110101100101;
		sqrt_table[ 146] = 36'b100110010000010001100110110101100010;
		sqrt_table[ 147] = 36'b100110010010111001011110110101011110;
		sqrt_table[ 148] = 36'b100110010101010010011000110101011011;
		sqrt_table[ 149] = 36'b100110010111111010111010110101010111;
		sqrt_table[ 150] = 36'b100110011010010100011110110101010100;
		sqrt_table[ 151] = 36'b100110011100111101101100110101010000;
		sqrt_table[ 152] = 36'b100110011111010111111010110101001101;
		sqrt_table[ 153] = 36'b100110100001110010010110110101001010;
		sqrt_table[ 154] = 36'b100110100100011100101000110101000110;
		sqrt_table[ 155] = 36'b100110100110110111101110110101000011;
		sqrt_table[ 156] = 36'b100110101001010011001000110100111111;
		sqrt_table[ 157] = 36'b100110101011101110111000110100111100;
		sqrt_table[ 158] = 36'b100110101110011010100000110100111000;
		sqrt_table[ 159] = 36'b100110110000100111001110110100110101;
		sqrt_table[ 160] = 36'b100110110011010011100110110100110010;
		sqrt_table[ 161] = 36'b100110110101110000100010110100101110;
		sqrt_table[ 162] = 36'b100110111000001101111000110100101011;
		sqrt_table[ 163] = 36'b100110111010101011011100110100101000;
		sqrt_table[ 164] = 36'b100110111101001001011000110100100100;
		sqrt_table[ 165] = 36'b100110111111100111100110110100100001;
		sqrt_table[ 166] = 36'b100111000010000110001010110100011110;
		sqrt_table[ 167] = 36'b100111000100010101000110110100011011;
		sqrt_table[ 168] = 36'b100111000111000100001100110100010111;
		sqrt_table[ 169] = 36'b100111001001010011101110110100010100;
		sqrt_table[ 170] = 36'b100111001100000011100000110100010000;
		sqrt_table[ 171] = 36'b100111001110010011100100110100001101;
		sqrt_table[ 172] = 36'b100111010000100011111110110100001010;
		sqrt_table[ 173] = 36'b100111010011010100110000110100000111;
		sqrt_table[ 174] = 36'b100111010101100101101100110100000100;
		sqrt_table[ 175] = 36'b100111011000000111000100110100000000;
		sqrt_table[ 176] = 36'b100111011010101000101110110011111101;
		sqrt_table[ 177] = 36'b100111011100111010100000110011111010;
		sqrt_table[ 178] = 36'b100111011111011100110010110011110111;
		sqrt_table[ 179] = 36'b100111100001101111001000110011110100;
		sqrt_table[ 180] = 36'b100111100100010010000100110011110000;
		sqrt_table[ 181] = 36'b100111100110100100111100110011101101;
		sqrt_table[ 182] = 36'b100111101001001000100000110011101010;
		sqrt_table[ 183] = 36'b100111101011011100000000110011100111;
		sqrt_table[ 184] = 36'b100111101110000000001000110011100100;
		sqrt_table[ 185] = 36'b100111110000010100001010110011100001;
		sqrt_table[ 186] = 36'b100111110010111000111100110011011101;
		sqrt_table[ 187] = 36'b100111110101001101100010110011011010;
		sqrt_table[ 188] = 36'b100111110111100010011010110011010111;
		sqrt_table[ 189] = 36'b100111111001110111100100110011010100;
		sqrt_table[ 190] = 36'b100111111100011101101010110011010001;
		sqrt_table[ 191] = 36'b100111111110110011010110110011001110;
		sqrt_table[ 192] = 36'b101000000001001001011000110011001011;
		sqrt_table[ 193] = 36'b101000000011110000010100110011001000;
		sqrt_table[ 194] = 36'b101000000101110110001010110011000101;
		sqrt_table[ 195] = 36'b101000001000011101110010110011000010;
		sqrt_table[ 196] = 36'b101000001010110100111000110010111111;
		sqrt_table[ 197] = 36'b101000001101001100010100110010111100;
		sqrt_table[ 198] = 36'b101000001111100011111110110010111001;
		sqrt_table[ 199] = 36'b101000010001111011111110110010110110;
		sqrt_table[ 200] = 36'b101000010100010100001100110010110011;
		sqrt_table[ 201] = 36'b101000010110101100110000110010110000;
		sqrt_table[ 202] = 36'b101000011000110100100110110010101101;
		sqrt_table[ 203] = 36'b101000011011011110101010110010101010;
		sqrt_table[ 204] = 36'b101000011101111000000010110010100111;
		sqrt_table[ 205] = 36'b101000100000010001101100110010100100;
		sqrt_table[ 206] = 36'b101000100010011010100010110010100001;
		sqrt_table[ 207] = 36'b101000100101000101111010110010011110;
		sqrt_table[ 208] = 36'b101000100111001111010000110010011011;
		sqrt_table[ 209] = 36'b101000101001101001111110110010011000;
		sqrt_table[ 210] = 36'b101000101100000101000110110010010101;
		sqrt_table[ 211] = 36'b101000101110001111001010110010010010;
		sqrt_table[ 212] = 36'b101000110000111100000100110010001111;
		sqrt_table[ 213] = 36'b101000110011000110101000110010001100;
		sqrt_table[ 214] = 36'b101000110101010001011110110010001010;
		sqrt_table[ 215] = 36'b101000110111111111010110110010000110;
		sqrt_table[ 216] = 36'b101000111001111001010000110010000100;
		sqrt_table[ 217] = 36'b101000111100100111101110110010000001;
		sqrt_table[ 218] = 36'b101000111110110011100100110001111110;
		sqrt_table[ 219] = 36'b101001000001010001001100110001111011;
		sqrt_table[ 220] = 36'b101001000011011101100000110001111000;
		sqrt_table[ 221] = 36'b101001000101111011101000110001110101;
		sqrt_table[ 222] = 36'b101001001000001000011110110001110011;
		sqrt_table[ 223] = 36'b101001001010010101100100110001110000;
		sqrt_table[ 224] = 36'b101001001100110100100110110001101101;
		sqrt_table[ 225] = 36'b101001001111010011110100110001101010;
		sqrt_table[ 226] = 36'b101001010001100001101010110001100111;
		sqrt_table[ 227] = 36'b101001010011101111110000110001100101;
		sqrt_table[ 228] = 36'b101001010110001111111010110001100010;
		sqrt_table[ 229] = 36'b101001011000011110100000110001011111;
		sqrt_table[ 230] = 36'b101001011010101101010100110001011100;
		sqrt_table[ 231] = 36'b101001011101001110010000110001011001;
		sqrt_table[ 232] = 36'b101001011111001011101100110001010111;
		sqrt_table[ 233] = 36'b101001100001111111001100110001010100;
		sqrt_table[ 234] = 36'b101001100011111101000000110001010001;
		sqrt_table[ 235] = 36'b101001100110001101000100110001001111;
		sqrt_table[ 236] = 36'b101001101000101111100000110001001100;
		sqrt_table[ 237] = 36'b101001101011000000000110110001001001;
		sqrt_table[ 238] = 36'b101001101101010000111010110001000110;
		sqrt_table[ 239] = 36'b101001101111100010000000110001000100;
		sqrt_table[ 240] = 36'b101001110001110011010110110001000001;
		sqrt_table[ 241] = 36'b101001110100010111000100110000111110;
		sqrt_table[ 242] = 36'b101001110110010110101100110000111100;
		sqrt_table[ 243] = 36'b101001111000101000110010110000111001;
		sqrt_table[ 244] = 36'b101001111011001101011010110000110110;
		sqrt_table[ 245] = 36'b101001111101001101101100110000110100;
		sqrt_table[ 246] = 36'b101001111111110010110110110000110001;
		sqrt_table[ 247] = 36'b101010000001110011100010110000101110;
		sqrt_table[ 248] = 36'b101010000100000110111000110000101100;
		sqrt_table[ 249] = 36'b101010000110011010011110110000101001;
		sqrt_table[ 250] = 36'b101010001001000000110010110000100110;
		sqrt_table[ 251] = 36'b101010001011000010011000110000100100;
		sqrt_table[ 252] = 36'b101010001101000100001000110000100001;
		sqrt_table[ 253] = 36'b101010001111101011010010110000011110;
		sqrt_table[ 254] = 36'b101010010001101101100000110000011100;
		sqrt_table[ 255] = 36'b101010010100010101010010110000011001;
		sqrt_table[ 256] = 36'b101010010110010111111010110000010111;
		sqrt_table[ 257] = 36'b101010011000101101100000110000010100;
		sqrt_table[ 258] = 36'b101010011010110000100110110000010010;
		sqrt_table[ 259] = 36'b101010011101000110101100110000001111;
		sqrt_table[ 260] = 36'b101010011111011101000000110000001100;
		sqrt_table[ 261] = 36'b101010100001110011100110110000001010;
		sqrt_table[ 262] = 36'b101010100011110111100010110000000111;
		sqrt_table[ 263] = 36'b101010100110001110101010110000000101;
		sqrt_table[ 264] = 36'b101010101000100110000000110000000010;
		sqrt_table[ 265] = 36'b101010101010101010101000110000000000;
		sqrt_table[ 266] = 36'b101010101100101111011100101111111101;
		sqrt_table[ 267] = 36'b101010101111011010100110101111111010;
		sqrt_table[ 268] = 36'b101010110001011111111000101111111000;
		sqrt_table[ 269] = 36'b101010110011100101011010101111110110;
		sqrt_table[ 270] = 36'b101010110101111110010000101111110011;
		sqrt_table[ 271] = 36'b101010111000000100001010101111110001;
		sqrt_table[ 272] = 36'b101010111010011101011110101111101110;
		sqrt_table[ 273] = 36'b101010111100100011111000101111101100;
		sqrt_table[ 274] = 36'b101010111110111101101110101111101001;
		sqrt_table[ 275] = 36'b101011000001000100100000101111100111;
		sqrt_table[ 276] = 36'b101011000011011110111000101111100100;
		sqrt_table[ 277] = 36'b101011000101100110001010101111100010;
		sqrt_table[ 278] = 36'b101011000111101101100110101111011111;
		sqrt_table[ 279] = 36'b101011001010001000101100101111011101;
		sqrt_table[ 280] = 36'b101011001100010000100110101111011010;
		sqrt_table[ 281] = 36'b101011001110011000110000101111011000;
		sqrt_table[ 282] = 36'b101011010000100001000110101111010110;
		sqrt_table[ 283] = 36'b101011010010111101001100101111010011;
		sqrt_table[ 284] = 36'b101011010101000101111100101111010001;
		sqrt_table[ 285] = 36'b101011010111100010100100101111001110;
		sqrt_table[ 286] = 36'b101011011001011000001100101111001100;
		sqrt_table[ 287] = 36'b101011011011110101001110101111001001;
		sqrt_table[ 288] = 36'b101011011101111110111100101111000111;
		sqrt_table[ 289] = 36'b101011100000001000110010101111000101;
		sqrt_table[ 290] = 36'b101011100010100110101010101111000010;
		sqrt_table[ 291] = 36'b101011100100011101001110101111000000;
		sqrt_table[ 292] = 36'b101011100110111011100010101110111101;
		sqrt_table[ 293] = 36'b101011101000110010011110101110111011;
		sqrt_table[ 294] = 36'b101011101011010001010100101110111001;
		sqrt_table[ 295] = 36'b101011101101011100100010101110110110;
		sqrt_table[ 296] = 36'b101011101111100111111100101110110100;
		sqrt_table[ 297] = 36'b101011110001110011100110101110110010;
		sqrt_table[ 298] = 36'b101011110011111111011010101110101111;
		sqrt_table[ 299] = 36'b101011110101110111011110101110101101;
		sqrt_table[ 300] = 36'b101011111000010111110010101110101011;
		sqrt_table[ 301] = 36'b101011111010100100010100101110101000;
		sqrt_table[ 302] = 36'b101011111100110001000010101110100110;
		sqrt_table[ 303] = 36'b101011111110111110000000101110100100;
		sqrt_table[ 304] = 36'b101100000001001011001000101110100001;
		sqrt_table[ 305] = 36'b101100000011000100010100101110011111;
		sqrt_table[ 306] = 36'b101100000101100110001100101110011101;
		sqrt_table[ 307] = 36'b101100000111011111110000101110011011;
		sqrt_table[ 308] = 36'b101100001010000010000100101110011000;
		sqrt_table[ 309] = 36'b101100001011111100000010101110010110;
		sqrt_table[ 310] = 36'b101100001110001010100000101110010100;
		sqrt_table[ 311] = 36'b101100010000000100110110101110010010;
		sqrt_table[ 312] = 36'b101100010010101000001100101110001111;
		sqrt_table[ 313] = 36'b101100010100100010110110101110001101;
		sqrt_table[ 314] = 36'b101100010110110010001010101110001011;
		sqrt_table[ 315] = 36'b101100011001000001110000101110001000;
		sqrt_table[ 316] = 36'b101100011011010001100010101110000110;
		sqrt_table[ 317] = 36'b101100011101001100111110101110000100;
		sqrt_table[ 318] = 36'b101100011111011101001110101110000010;
		sqrt_table[ 319] = 36'b101100100001101101101000101101111111;
		sqrt_table[ 320] = 36'b101100100011101001101000101101111101;
		sqrt_table[ 321] = 36'b101100100101111010100100101101111011;
		sqrt_table[ 322] = 36'b101100101000001011101000101101111001;
		sqrt_table[ 323] = 36'b101100101010001000001100101101110111;
		sqrt_table[ 324] = 36'b101100101100011001110000101101110100;
		sqrt_table[ 325] = 36'b101100101110101011100000101101110010;
		sqrt_table[ 326] = 36'b101100110000101000101010101101110000;
		sqrt_table[ 327] = 36'b101100110010100101111100101101101110;
		sqrt_table[ 328] = 36'b101100110101001101010010101101101011;
		sqrt_table[ 329] = 36'b101100110110110110000010101101101010;
		sqrt_table[ 330] = 36'b101100111001011101111000101101100111;
		sqrt_table[ 331] = 36'b101100111011011011111110101101100101;
		sqrt_table[ 332] = 36'b101100111101011010001100101101100011;
		sqrt_table[ 333] = 36'b101100111111101101101100101101100001;
		sqrt_table[ 334] = 36'b101101000001101100010100101101011111;
		sqrt_table[ 335] = 36'b101101000100000000010000101101011100;
		sqrt_table[ 336] = 36'b101101000101111111010010101101011010;
		sqrt_table[ 337] = 36'b101101000111111110011100101101011000;
		sqrt_table[ 338] = 36'b101101001010010011000010101101010110;
		sqrt_table[ 339] = 36'b101101001100100111111000101101010100;
		sqrt_table[ 340] = 36'b101101001110010010010110101101010010;
		sqrt_table[ 341] = 36'b101101010000111100111000101101001111;
		sqrt_table[ 342] = 36'b101101010010100111101110101101001110;
		sqrt_table[ 343] = 36'b101101010100111101011000101101001011;
		sqrt_table[ 344] = 36'b101101010110111101111000101101001001;
		sqrt_table[ 345] = 36'b101101011001010100000100101101000111;
		sqrt_table[ 346] = 36'b101101011010111111011000101101000101;
		sqrt_table[ 347] = 36'b101101011101010110000000101101000011;
		sqrt_table[ 348] = 36'b101101011111101100110000101101000001;
		sqrt_table[ 349] = 36'b101101100001011000101100101100111111;
		sqrt_table[ 350] = 36'b101101100011101111111000101100111101;
		sqrt_table[ 351] = 36'b101101100101110001101100101100111011;
		sqrt_table[ 352] = 36'b101101100111110011101100101100111001;
		sqrt_table[ 353] = 36'b101101101010001011100110101100110110;
		sqrt_table[ 354] = 36'b101101101100001101111100101100110100;
		sqrt_table[ 355] = 36'b101101101101111010110000101100110011;
		sqrt_table[ 356] = 36'b101101110000010011010010101100110000;
		sqrt_table[ 357] = 36'b101101110010101100000100101100101110;
		sqrt_table[ 358] = 36'b101101110100011001010100101100101100;
		sqrt_table[ 359] = 36'b101101110110011100101010101100101010;
		sqrt_table[ 360] = 36'b101101111000110110000100101100101000;
		sqrt_table[ 361] = 36'b101101111010100011110010101100100110;
		sqrt_table[ 362] = 36'b101101111100111101101000101100100100;
		sqrt_table[ 363] = 36'b101101111111000001101100101100100010;
		sqrt_table[ 364] = 36'b101110000001000101111100101100100000;
		sqrt_table[ 365] = 36'b101110000011001010011000101100011110;
		sqrt_table[ 366] = 36'b101110000101001111000010101100011100;
		sqrt_table[ 367] = 36'b101110000111010011110110101100011010;
		sqrt_table[ 368] = 36'b101110001001011000110110101100011000;
		sqrt_table[ 369] = 36'b101110001011011110000010101100010110;
		sqrt_table[ 370] = 36'b101110001101100011011010101100010100;
		sqrt_table[ 371] = 36'b101110001111010010101110101100010010;
		sqrt_table[ 372] = 36'b101110010001101110110000101100010000;
		sqrt_table[ 373] = 36'b101110010011110100101100101100001110;
		sqrt_table[ 374] = 36'b101110010101111010110100101100001100;
		sqrt_table[ 375] = 36'b101110011000000001001000101100001010;
		sqrt_table[ 376] = 36'b101110011001110001001100101100001000;
		sqrt_table[ 377] = 36'b101110011100001110010100101100000110;
		sqrt_table[ 378] = 36'b101110011101111110110000101100000100;
		sqrt_table[ 379] = 36'b101110100000000101110010101100000010;
		sqrt_table[ 380] = 36'b101110100010001101000100101100000000;
		sqrt_table[ 381] = 36'b101110100100010100011110101011111110;
		sqrt_table[ 382] = 36'b101110100110011100001000101011111100;
		sqrt_table[ 383] = 36'b101110101000100011111010101011111010;
		sqrt_table[ 384] = 36'b101110101010010101010000101011111001;
		sqrt_table[ 385] = 36'b101110101100011101011100101011110111;
		sqrt_table[ 386] = 36'b101110101110100101110100101011110101;
		sqrt_table[ 387] = 36'b101110110000101110011000101011110011;
		sqrt_table[ 388] = 36'b101110110010100000010110101011110001;
		sqrt_table[ 389] = 36'b101110110101000000000100101011101111;
		sqrt_table[ 390] = 36'b101110110110110010011010101011101101;
		sqrt_table[ 391] = 36'b101110111000111011101100101011101011;
		sqrt_table[ 392] = 36'b101110111010101110010000101011101001;
		sqrt_table[ 393] = 36'b101110111100110111111100101011100111;
		sqrt_table[ 394] = 36'b101110111111000001110100101011100101;
		sqrt_table[ 395] = 36'b101111000001001011111000101011100011;
		sqrt_table[ 396] = 36'b101111000010111111000110101011100010;
		sqrt_table[ 397] = 36'b101111000101001001100100101011100000;
		sqrt_table[ 398] = 36'b101111000110111101000010101011011110;
		sqrt_table[ 399] = 36'b101111001001000111110110101011011100;
		sqrt_table[ 400] = 36'b101111001011010010110110101011011010;
		sqrt_table[ 401] = 36'b101111001101000110110110101011011000;
		sqrt_table[ 402] = 36'b101111001111010010001110101011010110;
		sqrt_table[ 403] = 36'b101111010001011101110010101011010100;
		sqrt_table[ 404] = 36'b101111010011010010001110101011010011;
		sqrt_table[ 405] = 36'b101111010101011110001010101011010001;
		sqrt_table[ 406] = 36'b101111010111010011000000101011001111;
		sqrt_table[ 407] = 36'b101111011001011111010010101011001101;
		sqrt_table[ 408] = 36'b101111011011010100010110101011001011;
		sqrt_table[ 409] = 36'b101111011101100001000010101011001001;
		sqrt_table[ 410] = 36'b101111011111101101111010101011000111;
		sqrt_table[ 411] = 36'b101111100001100011011110101011000110;
		sqrt_table[ 412] = 36'b101111100011011001001100101011000100;
		sqrt_table[ 413] = 36'b101111100101100110101000101011000010;
		sqrt_table[ 414] = 36'b101111100111011100101000101011000000;
		sqrt_table[ 415] = 36'b101111101001101010011110101010111110;
		sqrt_table[ 416] = 36'b101111101011100000110000101010111101;
		sqrt_table[ 417] = 36'b101111101101101110111100101010111011;
		sqrt_table[ 418] = 36'b101111101111100101101010101010111001;
		sqrt_table[ 419] = 36'b101111110001011100011000101010110111;
		sqrt_table[ 420] = 36'b101111110011101011001000101010110101;
		sqrt_table[ 421] = 36'b101111110101111010000100101010110011;
		sqrt_table[ 422] = 36'b101111110111011001100010101010110010;
		sqrt_table[ 423] = 36'b101111111001101000110110101010110000;
		sqrt_table[ 424] = 36'b101111111011111000010110101010101110;
		sqrt_table[ 425] = 36'b101111111101110000000100101010101100;
		sqrt_table[ 426] = 36'b101111111111100111111110101010101011;
		sqrt_table[ 427] = 36'b110000000001100000000010101010101001;
		sqrt_table[ 428] = 36'b110000000011110000010100101010100111;
		sqrt_table[ 429] = 36'b110000000101101000100110101010100101;
		sqrt_table[ 430] = 36'b110000000111100001001100101010100100;
		sqrt_table[ 431] = 36'b110000001001110001111110101010100010;
		sqrt_table[ 432] = 36'b110000001011101010110100101010100000;
		sqrt_table[ 433] = 36'b110000001101100011110010101010011110;
		sqrt_table[ 434] = 36'b110000001111110101001100101010011100;
		sqrt_table[ 435] = 36'b110000010001010110010000101010011011;
		sqrt_table[ 436] = 36'b110000010011100111111110101010011001;
		sqrt_table[ 437] = 36'b110000010101100001100100101010010111;
		sqrt_table[ 438] = 36'b110000010111110011101100101010010101;
		sqrt_table[ 439] = 36'b110000011001010101001110101010010100;
		sqrt_table[ 440] = 36'b110000011011100111101110101010010010;
		sqrt_table[ 441] = 36'b110000011101100010000000101010010000;
		sqrt_table[ 442] = 36'b110000011111011100010110101010001111;
		sqrt_table[ 443] = 36'b110000100001101111011010101010001101;
		sqrt_table[ 444] = 36'b110000100011010001100110101010001011;
		sqrt_table[ 445] = 36'b110000100101100101000010101010001001;
		sqrt_table[ 446] = 36'b110000100111000111011100101010001000;
		sqrt_table[ 447] = 36'b110000101001011011010000101010000110;
		sqrt_table[ 448] = 36'b110000101011010110100110101010000100;
		sqrt_table[ 449] = 36'b110000101101101010110010101010000010;
		sqrt_table[ 450] = 36'b110000101111001101101110101010000001;
		sqrt_table[ 451] = 36'b110000110001001001100000101001111111;
		sqrt_table[ 452] = 36'b110000110011000101011110101001111110;
		sqrt_table[ 453] = 36'b110000110101011010011010101001111100;
		sqrt_table[ 454] = 36'b110000110110111101110100101001111010;
		sqrt_table[ 455] = 36'b110000111001010011001000101001111000;
		sqrt_table[ 456] = 36'b110000111011001111101110101001110111;
		sqrt_table[ 457] = 36'b110000111100110011011110101001110101;
		sqrt_table[ 458] = 36'b110000111111001001010110101001110011;
		sqrt_table[ 459] = 36'b110001000001000110011110101001110010;
		sqrt_table[ 460] = 36'b110001000010101010101000101001110000;
		sqrt_table[ 461] = 36'b110001000101000001000010101001101110;
		sqrt_table[ 462] = 36'b110001000110111110100100101001101101;
		sqrt_table[ 463] = 36'b110001001000100011000100101001101011;
		sqrt_table[ 464] = 36'b110001001010111010000100101001101001;
		sqrt_table[ 465] = 36'b110001001100111000001000101001101000;
		sqrt_table[ 466] = 36'b110001001110011101000010101001100110;
		sqrt_table[ 467] = 36'b110001010000110100100100101001100100;
		sqrt_table[ 468] = 36'b110001010010011001110000101001100011;
		sqrt_table[ 469] = 36'b110001010100011000010110101001100001;
		sqrt_table[ 470] = 36'b110001010110010111001000101001100000;
		sqrt_table[ 471] = 36'b110001011000101111011110101001011110;
		sqrt_table[ 472] = 36'b110001011010010101001000101001011100;
		sqrt_table[ 473] = 36'b110001011100010100010110101001011011;
		sqrt_table[ 474] = 36'b110001011101111010010000101001011001;
		sqrt_table[ 475] = 36'b110001100000010011010100101001010111;
		sqrt_table[ 476] = 36'b110001100001111001011110101001010110;
		sqrt_table[ 477] = 36'b110001100100010010111010101001010100;
		sqrt_table[ 478] = 36'b110001100101111001010110101001010011;
		sqrt_table[ 479] = 36'b110001100111111001100010101001010001;
		sqrt_table[ 480] = 36'b110001101001111001110110101001001111;
		sqrt_table[ 481] = 36'b110001101011111010010110101001001110;
		sqrt_table[ 482] = 36'b110001101101100001010000101001001100;
		sqrt_table[ 483] = 36'b110001101111100010000100101001001011;
		sqrt_table[ 484] = 36'b110001110001100011000010101001001001;
		sqrt_table[ 485] = 36'b110001110011100100001000101001000111;
		sqrt_table[ 486] = 36'b110001110101100101011010101001000110;
		sqrt_table[ 487] = 36'b110001110111001100111100101001000100;
		sqrt_table[ 488] = 36'b110001111001001110100010101001000011;
		sqrt_table[ 489] = 36'b110001111011010000010010101001000001;
		sqrt_table[ 490] = 36'b110001111101010010001010101000111111;
		sqrt_table[ 491] = 36'b110001111110111010001100101000111110;
		sqrt_table[ 492] = 36'b110010000000111100011100101000111100;
		sqrt_table[ 493] = 36'b110010000010111110110000101000111011;
		sqrt_table[ 494] = 36'b110010000100100111001100101000111001;
		sqrt_table[ 495] = 36'b110010000110101001111000101000111000;
		sqrt_table[ 496] = 36'b110010001000101100101110101000110110;
		sqrt_table[ 497] = 36'b110010001010101111101100101000110100;
		sqrt_table[ 498] = 36'b110010001100011000101000101000110011;
		sqrt_table[ 499] = 36'b110010001110011011111010101000110001;
		sqrt_table[ 500] = 36'b110010010000000101000100101000110000;
		sqrt_table[ 501] = 36'b110010010010001000101100101000101110;
		sqrt_table[ 502] = 36'b110010010100001100011100101000101101;
		sqrt_table[ 503] = 36'b110010010101110110000000101000101011;
		sqrt_table[ 504] = 36'b110010010111111010000110101000101010;
		sqrt_table[ 505] = 36'b110010011001111110010110101000101000;
		sqrt_table[ 506] = 36'b110010011011101000001110101000100111;
		sqrt_table[ 507] = 36'b110010011101101100110100101000100101;
		sqrt_table[ 508] = 36'b110010011111110001011110101000100011;
		sqrt_table[ 509] = 36'b110010100001011011110100101000100010;
		sqrt_table[ 510] = 36'b110010100011000110001100101000100001;
		sqrt_table[ 511] = 36'b110010100101001011011010101000011111;
		sqrt_table[ 512] = 36'b110010100111010000101100101000011101;
		sqrt_table[ 513] = 36'b110010101000111011100010101000011100;
		sqrt_table[ 514] = 36'b110010101011000001001010101000011010;
		sqrt_table[ 515] = 36'b110010101100101100001110101000011001;
		sqrt_table[ 516] = 36'b110010101110110010001010101000010111;
		sqrt_table[ 517] = 36'b110010110000011101011100101000010110;
		sqrt_table[ 518] = 36'b110010110010100011101110101000010100;
		sqrt_table[ 519] = 36'b110010110100001111010010101000010011;
		sqrt_table[ 520] = 36'b110010110110010101110100101000010001;
		sqrt_table[ 521] = 36'b110010111000000001101010101000010000;
		sqrt_table[ 522] = 36'b110010111010001000100010101000001110;
		sqrt_table[ 523] = 36'b110010111011110100100110101000001101;
		sqrt_table[ 524] = 36'b110010111101111011110010101000001011;
		sqrt_table[ 525] = 36'b110010111111101000000100101000001010;
		sqrt_table[ 526] = 36'b110011000001101111101000101000001000;
		sqrt_table[ 527] = 36'b110011000011011100001100101000000111;
		sqrt_table[ 528] = 36'b110011000101001000110110101000000110;
		sqrt_table[ 529] = 36'b110011000111010000110010101000000100;
		sqrt_table[ 530] = 36'b110011001000111101101110101000000011;
		sqrt_table[ 531] = 36'b110011001011000110000010101000000001;
		sqrt_table[ 532] = 36'b110011001100110011001100101000000000;
		sqrt_table[ 533] = 36'b110011001110111011110100100111111110;
		sqrt_table[ 534] = 36'b110011010000101001001100100111111101;
		sqrt_table[ 535] = 36'b110011010010010110110000100111111011;
		sqrt_table[ 536] = 36'b110011010100000100011010100111111010;
		sqrt_table[ 537] = 36'b110011010110001101101010100111111000;
		sqrt_table[ 538] = 36'b110011011000010111000010100111110111;
		sqrt_table[ 539] = 36'b110011011001101001100110100111110110;
		sqrt_table[ 540] = 36'b110011011011110011010100100111110100;
		sqrt_table[ 541] = 36'b110011011101111101001010100111110010;
		sqrt_table[ 542] = 36'b110011011111001111111100100111110001;
		sqrt_table[ 543] = 36'b110011100001011010001010100111110000;
		sqrt_table[ 544] = 36'b110011100011100100011110100111101110;
		sqrt_table[ 545] = 36'b110011100100110111100110100111101101;
		sqrt_table[ 546] = 36'b110011100111000010001110100111101011;
		sqrt_table[ 547] = 36'b110011101000110001010000100111101010;
		sqrt_table[ 548] = 36'b110011101010111100010000100111101000;
		sqrt_table[ 549] = 36'b110011101100001111101100100111100111;
		sqrt_table[ 550] = 36'b110011101110011010111110100111100110;
		sqrt_table[ 551] = 36'b110011110000100110011010100111100100;
		sqrt_table[ 552] = 36'b110011110001111010001100100111100011;
		sqrt_table[ 553] = 36'b110011110100000101110110100111100001;
		sqrt_table[ 554] = 36'b110011110101110101110100100111100000;
		sqrt_table[ 555] = 36'b110011110111100101110100100111011111;
		sqrt_table[ 556] = 36'b110011111001010110000000100111011101;
		sqrt_table[ 557] = 36'b110011111011100010011000100111011100;
		sqrt_table[ 558] = 36'b110011111101010010110010100111011010;
		sqrt_table[ 559] = 36'b110011111111000011010110100111011001;
		sqrt_table[ 560] = 36'b110100000000110100000000100111011000;
		sqrt_table[ 561] = 36'b110100000011000001000000100111010110;
		sqrt_table[ 562] = 36'b110100000100010101101110100111010101;
		sqrt_table[ 563] = 36'b110100000110100010111100100111010011;
		sqrt_table[ 564] = 36'b110100001000010100001010100111010010;
		sqrt_table[ 565] = 36'b110100001010000101011010100111010001;
		sqrt_table[ 566] = 36'b110100001011110110110110100111001111;
		sqrt_table[ 567] = 36'b110100001110000100110010100111001110;
		sqrt_table[ 568] = 36'b110100001111011010000000100111001101;
		sqrt_table[ 569] = 36'b110100010001101000010010100111001011;
		sqrt_table[ 570] = 36'b110100010011011010001100100111001010;
		sqrt_table[ 571] = 36'b110100010101001100010000100111001000;
		sqrt_table[ 572] = 36'b110100010110111110011100100111000111;
		sqrt_table[ 573] = 36'b110100011000110000101110100111000110;
		sqrt_table[ 574] = 36'b110100011010100011000110100111000100;
		sqrt_table[ 575] = 36'b110100011100110010010000100111000011;
		sqrt_table[ 576] = 36'b110100011110001000010010100111000010;
		sqrt_table[ 577] = 36'b110100100000010111110010100111000000;
		sqrt_table[ 578] = 36'b110100100001101110000000100110111111;
		sqrt_table[ 579] = 36'b110100100011111101101110100110111101;
		sqrt_table[ 580] = 36'b110100100101110000111100100110111100;
		sqrt_table[ 581] = 36'b110100100111000111011100100110111011;
		sqrt_table[ 582] = 36'b110100101001010111101000100110111001;
		sqrt_table[ 583] = 36'b110100101011001011001110100110111000;
		sqrt_table[ 584] = 36'b110100101100111110110110100110110111;
		sqrt_table[ 585] = 36'b110100101110110010101010100110110101;
		sqrt_table[ 586] = 36'b110100110000100110100100100110110100;
		sqrt_table[ 587] = 36'b110100110010011010101000100110110011;
		sqrt_table[ 588] = 36'b110100110100001110110000100110110001;
		sqrt_table[ 589] = 36'b110100110110000011000110100110110000;
		sqrt_table[ 590] = 36'b110100110111011010011100100110101111;
		sqrt_table[ 591] = 36'b110100111001101100000010100110101101;
		sqrt_table[ 592] = 36'b110100111011100000110000100110101100;
		sqrt_table[ 593] = 36'b110100111101010101100000100110101011;
		sqrt_table[ 594] = 36'b110100111111001010011100100110101001;
		sqrt_table[ 595] = 36'b110101000000111111011110100110101000;
		sqrt_table[ 596] = 36'b110101000010110100101010100110100111;
		sqrt_table[ 597] = 36'b110101000100001100101010100110100110;
		sqrt_table[ 598] = 36'b110101000110011111011000100110100100;
		sqrt_table[ 599] = 36'b110101001000010100111100100110100011;
		sqrt_table[ 600] = 36'b110101001001101101001110100110100010;
		sqrt_table[ 601] = 36'b110101001100000000011010100110100000;
		sqrt_table[ 602] = 36'b110101001101011000111000100110011111;
		sqrt_table[ 603] = 36'b110101001111001110111010100110011110;
		sqrt_table[ 604] = 36'b110101010001000101000100100110011100;
		sqrt_table[ 605] = 36'b110101010010111011011000100110011011;
		sqrt_table[ 606] = 36'b110101010100110001110010100110011010;
		sqrt_table[ 607] = 36'b110101010110101000010100100110011000;
		sqrt_table[ 608] = 36'b110101011000011111000000100110010111;
		sqrt_table[ 609] = 36'b110101011010010101110010100110010110;
		sqrt_table[ 610] = 36'b110101011011101110111100100110010101;
		sqrt_table[ 611] = 36'b110101011101100110000000100110010011;
		sqrt_table[ 612] = 36'b110101011111111010111110100110010010;
		sqrt_table[ 613] = 36'b110101100001010100011010100110010001;
		sqrt_table[ 614] = 36'b110101100011001011110110100110001111;
		sqrt_table[ 615] = 36'b110101100100100101100000100110001110;
		sqrt_table[ 616] = 36'b110101100110111011000100100110001101;
		sqrt_table[ 617] = 36'b110101101000010100111100100110001100;
		sqrt_table[ 618] = 36'b110101101010101010110110100110001010;
		sqrt_table[ 619] = 36'b110101101100000100111010100110001001;
		sqrt_table[ 620] = 36'b110101101101011111000000100110001000;
		sqrt_table[ 621] = 36'b110101101111110101010110100110000110;
		sqrt_table[ 622] = 36'b110101110001001111101000100110000101;
		sqrt_table[ 623] = 36'b110101110011100110010110100110000100;
		sqrt_table[ 624] = 36'b110101110101000000110110100110000011;
		sqrt_table[ 625] = 36'b110101110110111001100110100110000001;
		sqrt_table[ 626] = 36'b110101111000010100010100100110000000;
		sqrt_table[ 627] = 36'b110101111010001101011000100101111111;
		sqrt_table[ 628] = 36'b110101111100100100110100100101111101;
		sqrt_table[ 629] = 36'b110101111101100001011110100101111101;
		sqrt_table[ 630] = 36'b110101111111111001010000100101111011;
		sqrt_table[ 631] = 36'b110110000001010100011000100101111010;
		sqrt_table[ 632] = 36'b110110000011001110000100100101111001;
		sqrt_table[ 633] = 36'b110110000101000111110100100101110111;
		sqrt_table[ 634] = 36'b110110000111000001110010100101110110;
		sqrt_table[ 635] = 36'b110110001000011101010110100101110101;
		sqrt_table[ 636] = 36'b110110001010010111011110100101110100;
		sqrt_table[ 637] = 36'b110110001100010001110010100101110010;
		sqrt_table[ 638] = 36'b110110001101101101100100100101110001;
		sqrt_table[ 639] = 36'b110110001111101000000110100101110000;
		sqrt_table[ 640] = 36'b110110010001100010110010100101101111;
		sqrt_table[ 641] = 36'b110110010010111110111000100101101110;
		sqrt_table[ 642] = 36'b110110010101011000100000100101101100;
		sqrt_table[ 643] = 36'b110110010110010110000000100101101011;
		sqrt_table[ 644] = 36'b110110011000110000000000100101101010;
		sqrt_table[ 645] = 36'b110110011010001100011110100101101001;
		sqrt_table[ 646] = 36'b110110011100000111110110100101100111;
		sqrt_table[ 647] = 36'b110110011101100100100010100101100110;
		sqrt_table[ 648] = 36'b110110011111100000001110100101100101;
		sqrt_table[ 649] = 36'b110110100001011100000000100101100100;
		sqrt_table[ 650] = 36'b110110100011010111111010100101100010;
		sqrt_table[ 651] = 36'b110110100100110100111010100101100001;
		sqrt_table[ 652] = 36'b110110100110010010000100100101100000;
		sqrt_table[ 653] = 36'b110110101000001110011000100101011111;
		sqrt_table[ 654] = 36'b110110101010001010110010100101011110;
		sqrt_table[ 655] = 36'b110110101100000111010100100101011100;
		sqrt_table[ 656] = 36'b110110101101100100110010100101011011;
		sqrt_table[ 657] = 36'b110110101111100001101000100101011010;
		sqrt_table[ 658] = 36'b110110110000111111010110100101011001;
		sqrt_table[ 659] = 36'b110110110010111100011000100101011000;
		sqrt_table[ 660] = 36'b110110110100011010001110100101010111;
		sqrt_table[ 661] = 36'b110110110110010111011110100101010101;
		sqrt_table[ 662] = 36'b110110111000010100111100100101010100;
		sqrt_table[ 663] = 36'b110110111001110011000110100101010011;
		sqrt_table[ 664] = 36'b110110111011110000110000100101010010;
		sqrt_table[ 665] = 36'b110110111101001111000110100101010001;
		sqrt_table[ 666] = 36'b110110111111001100111110100101001111;
		sqrt_table[ 667] = 36'b110111000000101011100010100101001110;
		sqrt_table[ 668] = 36'b110111000010101001101110100101001101;
		sqrt_table[ 669] = 36'b110111000100101000000000100101001100;
		sqrt_table[ 670] = 36'b110111000110000110110010100101001011;
		sqrt_table[ 671] = 36'b110111000111100101101110100101001010;
		sqrt_table[ 672] = 36'b110111001001100100011000100101001000;
		sqrt_table[ 673] = 36'b110111001011100011001100100101000111;
		sqrt_table[ 674] = 36'b110111001101000010010110100101000110;
		sqrt_table[ 675] = 36'b110111001111000001011010100101000101;
		sqrt_table[ 676] = 36'b110111010000100000110100100101000100;
		sqrt_table[ 677] = 36'b110111010010000000010000100101000011;
		sqrt_table[ 678] = 36'b110111010011111111101000100101000001;
		sqrt_table[ 679] = 36'b110111010101111111001110100101000000;
		sqrt_table[ 680] = 36'b110111010111011111000000100100111111;
		sqrt_table[ 681] = 36'b110111011000111110110100100100111110;
		sqrt_table[ 682] = 36'b110111011010111110101100100100111101;
		sqrt_table[ 683] = 36'b110111011100111110110000100100111011;
		sqrt_table[ 684] = 36'b110111011101111110110110100100111011;
		sqrt_table[ 685] = 36'b110111100000011111001110100100111001;
		sqrt_table[ 686] = 36'b110111100001011111011010100100111000;
		sqrt_table[ 687] = 36'b110111100100000000000100100100110111;
		sqrt_table[ 688] = 36'b110111100101000000011010100100110110;
		sqrt_table[ 689] = 36'b110111100111000001001110100100110101;
		sqrt_table[ 690] = 36'b110111101001000010000110100100110011;
		sqrt_table[ 691] = 36'b110111101010100010111010100100110010;
		sqrt_table[ 692] = 36'b110111101100000011110000100100110001;
		sqrt_table[ 693] = 36'b110111101110000101000110100100110000;
		sqrt_table[ 694] = 36'b110111101111100110001010100100101111;
		sqrt_table[ 695] = 36'b110111110001100111101110100100101110;
		sqrt_table[ 696] = 36'b110111110011001000111100100100101101;
		sqrt_table[ 697] = 36'b110111110100101010010100100100101100;
		sqrt_table[ 698] = 36'b110111110110101100001110100100101010;
		sqrt_table[ 699] = 36'b110111111000001101101110100100101001;
		sqrt_table[ 700] = 36'b110111111001101111010110100100101000;
		sqrt_table[ 701] = 36'b110111111011110001101010100100100111;
		sqrt_table[ 702] = 36'b110111111101010011011110100100100110;
		sqrt_table[ 703] = 36'b110111111111010101111110100100100101;
		sqrt_table[ 704] = 36'b111000000000111000000000100100100100;
		sqrt_table[ 705] = 36'b111000000010011010000100100100100011;
		sqrt_table[ 706] = 36'b111000000100011101000000100100100001;
		sqrt_table[ 707] = 36'b111000000101111111010010100100100000;
		sqrt_table[ 708] = 36'b111000000111100001101010100100011111;
		sqrt_table[ 709] = 36'b111000001001100100111100100100011110;
		sqrt_table[ 710] = 36'b111000001011000111100010100100011101;
		sqrt_table[ 711] = 36'b111000001100101010001010100100011100;
		sqrt_table[ 712] = 36'b111000001110101101110110100100011011;
		sqrt_table[ 713] = 36'b111000010000010000101100100100011010;
		sqrt_table[ 714] = 36'b111000010001110011101000100100011001;
		sqrt_table[ 715] = 36'b111000010011110111101000100100010111;
		sqrt_table[ 716] = 36'b111000010101011010110010100100010110;
		sqrt_table[ 717] = 36'b111000010110111101111110100100010101;
		sqrt_table[ 718] = 36'b111000011000100001010100100100010100;
		sqrt_table[ 719] = 36'b111000011010100101111000100100010011;
		sqrt_table[ 720] = 36'b111000011100001001010110100100010010;
		sqrt_table[ 721] = 36'b111000011110001110001010100100010001;
		sqrt_table[ 722] = 36'b111000011111010000101000100100010000;
		sqrt_table[ 723] = 36'b111000100001010101101000100100001111;
		sqrt_table[ 724] = 36'b111000100010111001100010100100001110;
		sqrt_table[ 725] = 36'b111000100100111110110100100100001100;
		sqrt_table[ 726] = 36'b111000100110000001100010100100001100;
		sqrt_table[ 727] = 36'b111000101000000111000100100100001010;
		sqrt_table[ 728] = 36'b111000101001101011010100100100001001;
		sqrt_table[ 729] = 36'b111000101011110001000110100100001000;
		sqrt_table[ 730] = 36'b111000101100110100000010100100000111;
		sqrt_table[ 731] = 36'b111000101110111010001000100100000110;
		sqrt_table[ 732] = 36'b111000110000011110110000100100000101;
		sqrt_table[ 733] = 36'b111000110010100101000010100100000100;
		sqrt_table[ 734] = 36'b111000110011101000010000100100000011;
		sqrt_table[ 735] = 36'b111000110101101110110010100100000010;
		sqrt_table[ 736] = 36'b111000110111010011110000100100000001;
		sqrt_table[ 737] = 36'b111000111000111000111000100100000000;
		sqrt_table[ 738] = 36'b111000111010011110000010100011111111;
		sqrt_table[ 739] = 36'b111000111100100101000110100011111101;
		sqrt_table[ 740] = 36'b111000111110001010100000100011111100;
		sqrt_table[ 741] = 36'b111000111111101111111100100011111011;
		sqrt_table[ 742] = 36'b111001000001010101100010100011111010;
		sqrt_table[ 743] = 36'b111001000010111011001010100011111001;
		sqrt_table[ 744] = 36'b111001000101000010110100100011111000;
		sqrt_table[ 745] = 36'b111001000110000110101100100011110111;
		sqrt_table[ 746] = 36'b111001001000001110101010100011110110;
		sqrt_table[ 747] = 36'b111001001001110100101100100011110101;
		sqrt_table[ 748] = 36'b111001001011011010110100100011110100;
		sqrt_table[ 749] = 36'b111001001101000001000010100011110011;
		sqrt_table[ 750] = 36'b111001001111001001011100100011110010;
		sqrt_table[ 751] = 36'b111001010000001101101110100011110001;
		sqrt_table[ 752] = 36'b111001010010010110011000100011110000;
		sqrt_table[ 753] = 36'b111001010011111100111100100011101111;
		sqrt_table[ 754] = 36'b111001010101100011101010100011101110;
		sqrt_table[ 755] = 36'b111001010111001010011010100011101101;
		sqrt_table[ 756] = 36'b111001011000110001010100100011101100;
		sqrt_table[ 757] = 36'b111001011010111010100110100011101010;
		sqrt_table[ 758] = 36'b111001011011111111010100100011101010;
		sqrt_table[ 759] = 36'b111001011110001000110110100011101000;
		sqrt_table[ 760] = 36'b111001011111001101101100100011101000;
		sqrt_table[ 761] = 36'b111001100001010111011110100011100110;
		sqrt_table[ 762] = 36'b111001100010111110111000100011100101;
		sqrt_table[ 763] = 36'b111001100100100110011100100011100100;
		sqrt_table[ 764] = 36'b111001100110001110000010100011100011;
		sqrt_table[ 765] = 36'b111001100111110101110010100011100010;
		sqrt_table[ 766] = 36'b111001101010000000001110100011100001;
		sqrt_table[ 767] = 36'b111001101011000101100000100011100000;
		sqrt_table[ 768] = 36'b111001101100101101011110100011011111;
		sqrt_table[ 769] = 36'b111001101110111000010000100011011110;
		sqrt_table[ 770] = 36'b111001101111111101101100100011011101;
		sqrt_table[ 771] = 36'b111001110010001000110010100011011100;
		sqrt_table[ 772] = 36'b111001110011001110010110100011011011;
		sqrt_table[ 773] = 36'b111001110101011001101000100011011010;
		sqrt_table[ 774] = 36'b111001110111000010001110100011011001;
		sqrt_table[ 775] = 36'b111001111000101010110110100011011000;
		sqrt_table[ 776] = 36'b111001111001110000101010100011010111;
		sqrt_table[ 777] = 36'b111001111011111100100000100011010110;
		sqrt_table[ 778] = 36'b111001111101100101011100100011010101;
		sqrt_table[ 779] = 36'b111001111111001110011110100011010100;
		sqrt_table[ 780] = 36'b111010000000110111100110100011010011;
		sqrt_table[ 781] = 36'b111010000010100000110100100011010010;
		sqrt_table[ 782] = 36'b111010000100001010001010100011010001;
		sqrt_table[ 783] = 36'b111010000101110011100010100011010000;
		sqrt_table[ 784] = 36'b111010000111011101000100100011001111;
		sqrt_table[ 785] = 36'b111010001001000110101000100011001110;
		sqrt_table[ 786] = 36'b111010001010110000010110100011001101;
		sqrt_table[ 787] = 36'b111010001100011010000110100011001100;
		sqrt_table[ 788] = 36'b111010001110000100000000100011001011;
		sqrt_table[ 789] = 36'b111010001111101101111100100011001010;
		sqrt_table[ 790] = 36'b111010010001011000000010100011001001;
		sqrt_table[ 791] = 36'b111010010010011110110000100011001000;
		sqrt_table[ 792] = 36'b111010010100101100011100100011000111;
		sqrt_table[ 793] = 36'b111010010110010110110000100011000110;
		sqrt_table[ 794] = 36'b111010011000000001001110100011000101;
		sqrt_table[ 795] = 36'b111010011001101011101110100011000100;
		sqrt_table[ 796] = 36'b111010011011010110011000100011000011;
		sqrt_table[ 797] = 36'b111010011100011101100000100011000010;
		sqrt_table[ 798] = 36'b111010011110101011111100100011000001;
		sqrt_table[ 799] = 36'b111010100000010110110110100011000000;
		sqrt_table[ 800] = 36'b111010100001011110001010100010111111;
		sqrt_table[ 801] = 36'b111010100011101100111100100010111110;
		sqrt_table[ 802] = 36'b111010100100110100011000100010111101;
		sqrt_table[ 803] = 36'b111010100110011111101100100010111100;
		sqrt_table[ 804] = 36'b111010101000101110111000100010111011;
		sqrt_table[ 805] = 36'b111010101001110110100010100010111010;
		sqrt_table[ 806] = 36'b111010101011100010000100100010111001;
		sqrt_table[ 807] = 36'b111010101101001101101110100010111000;
		sqrt_table[ 808] = 36'b111010101110111001011110100010110111;
		sqrt_table[ 809] = 36'b111010110000100101010100100010110110;
		sqrt_table[ 810] = 36'b111010110010010001010000100010110101;
		sqrt_table[ 811] = 36'b111010110011011001010010100010110101;
		sqrt_table[ 812] = 36'b111010110101101001011010100010110011;
		sqrt_table[ 813] = 36'b111010110110110001100100100010110011;
		sqrt_table[ 814] = 36'b111010111001000010000000100010110001;
		sqrt_table[ 815] = 36'b111010111010001010010010100010110001;
		sqrt_table[ 816] = 36'b111010111011110110110010100010110000;
		sqrt_table[ 817] = 36'b111010111101100011011000100010101111;
		sqrt_table[ 818] = 36'b111010111111010000000100100010101110;
		sqrt_table[ 819] = 36'b111011000000111100110110100010101101;
		sqrt_table[ 820] = 36'b111011000010000101011100100010101100;
		sqrt_table[ 821] = 36'b111011000100010110101100100010101011;
		sqrt_table[ 822] = 36'b111011000101011111011010100010101010;
		sqrt_table[ 823] = 36'b111011000111001100100110100010101001;
		sqrt_table[ 824] = 36'b111011001000111001110100100010101000;
		sqrt_table[ 825] = 36'b111011001010100111001100100010100111;
		sqrt_table[ 826] = 36'b111011001100010100100110100010100110;
		sqrt_table[ 827] = 36'b111011001110000010001010100010100101;
		sqrt_table[ 828] = 36'b111011001111001011001110100010100100;
		sqrt_table[ 829] = 36'b111011010000111000111100100010100011;
		sqrt_table[ 830] = 36'b111011010011001011010110100010100010;
		sqrt_table[ 831] = 36'b111011010100010100100110100010100001;
		sqrt_table[ 832] = 36'b111011010101011101111100100010100001;
		sqrt_table[ 833] = 36'b111011010111110000110000100010011111;
		sqrt_table[ 834] = 36'b111011011000111010001110100010011111;
		sqrt_table[ 835] = 36'b111011011010101000100000100010011110;
		sqrt_table[ 836] = 36'b111011011100010110111000100010011101;
		sqrt_table[ 837] = 36'b111011011110000101010110100010011100;
		sqrt_table[ 838] = 36'b111011011111110011111010100010011011;
		sqrt_table[ 839] = 36'b111011100000111101101100100010011010;
		sqrt_table[ 840] = 36'b111011100011010001010100100010011001;
		sqrt_table[ 841] = 36'b111011100100011011001110100010011000;
		sqrt_table[ 842] = 36'b111011100101100101001010100010010111;
		sqrt_table[ 843] = 36'b111011100111111001010000100010010110;
		sqrt_table[ 844] = 36'b111011101001000011010100100010010101;
		sqrt_table[ 845] = 36'b111011101010110010100010100010010100;
		sqrt_table[ 846] = 36'b111011101100100001110110100010010011;
		sqrt_table[ 847] = 36'b111011101110010001010000100010010010;
		sqrt_table[ 848] = 36'b111011110000000000110000100010010001;
		sqrt_table[ 849] = 36'b111011110001001011001010100010010001;
		sqrt_table[ 850] = 36'b111011110010111010111000100010010000;
		sqrt_table[ 851] = 36'b111011110100101010101000100010001111;
		sqrt_table[ 852] = 36'b111011110101110101001110100010001110;
		sqrt_table[ 853] = 36'b111011110111100101001100100010001101;
		sqrt_table[ 854] = 36'b111011111001010101010000100010001100;
		sqrt_table[ 855] = 36'b111011111011000101011010100010001011;
		sqrt_table[ 856] = 36'b111011111100010000001110100010001010;
		sqrt_table[ 857] = 36'b111011111110100110000010100010001001;
		sqrt_table[ 858] = 36'b111011111111110001000000100010001000;
		sqrt_table[ 859] = 36'b111100000000111100000000100010001000;
		sqrt_table[ 860] = 36'b111100000011010010001010100010000110;
		sqrt_table[ 861] = 36'b111100000100011101010110100010000110;
		sqrt_table[ 862] = 36'b111100000110001110001000100010000101;
		sqrt_table[ 863] = 36'b111100000111011001011010100010000100;
		sqrt_table[ 864] = 36'b111100001001001010011010100010000011;
		sqrt_table[ 865] = 36'b111100001010111011100000100010000010;
		sqrt_table[ 866] = 36'b111100001100101100101100100010000001;
		sqrt_table[ 867] = 36'b111100001110011101111110100010000000;
		sqrt_table[ 868] = 36'b111100001111101001100010100001111111;
		sqrt_table[ 869] = 36'b111100010000110101001100100001111111;
		sqrt_table[ 870] = 36'b111100010011001100100100100001111101;
		sqrt_table[ 871] = 36'b111100010100011000010110100001111101;
		sqrt_table[ 872] = 36'b111100010110001010001000100001111100;
		sqrt_table[ 873] = 36'b111100010111010110000010100001111011;
		sqrt_table[ 874] = 36'b111100011001101101111100100001111010;
		sqrt_table[ 875] = 36'b111100011010111001111110100001111001;
		sqrt_table[ 876] = 36'b111100011100000110000100100001111000;
		sqrt_table[ 877] = 36'b111100011101111000010000100001110111;
		sqrt_table[ 878] = 36'b111100011111101010100100100001110110;
		sqrt_table[ 879] = 36'b111100100001011100111110100001110101;
		sqrt_table[ 880] = 36'b111100100010101001010100100001110101;
		sqrt_table[ 881] = 36'b111100100100011011111010100001110100;
		sqrt_table[ 882] = 36'b111100100101101000011000100001110011;
		sqrt_table[ 883] = 36'b111100101000000001011010100001110010;
		sqrt_table[ 884] = 36'b111100101000100111101100100001110001;
		sqrt_table[ 885] = 36'b111100101011000000111110100001110000;
		sqrt_table[ 886] = 36'b111100101100001101101010100001101111;
		sqrt_table[ 887] = 36'b111100101110000000110110100001101110;
		sqrt_table[ 888] = 36'b111100101111001101101100100001101110;
		sqrt_table[ 889] = 36'b111100110001000001000010100001101101;
		sqrt_table[ 890] = 36'b111100110010110100011110100001101100;
		sqrt_table[ 891] = 36'b111100110100000001100000100001101011;
		sqrt_table[ 892] = 36'b111100110101110101000110100001101010;
		sqrt_table[ 893] = 36'b111100110111000010001110100001101001;
		sqrt_table[ 894] = 36'b111100111000110110000100100001101000;
		sqrt_table[ 895] = 36'b111100111010101001111100100001100111;
		sqrt_table[ 896] = 36'b111100111100011101111110100001100110;
		sqrt_table[ 897] = 36'b111100111101000100101100100001100110;
		sqrt_table[ 898] = 36'b111100111111011111100100100001100101;
		sqrt_table[ 899] = 36'b111101000000101101000110100001100100;
		sqrt_table[ 900] = 36'b111101000010100001100000100001100011;
		sqrt_table[ 901] = 36'b111101000011101111001000100001100010;
		sqrt_table[ 902] = 36'b111101000101100011101100100001100001;
		sqrt_table[ 903] = 36'b111101000111011000010110100001100000;
		sqrt_table[ 904] = 36'b111101001000100110001100100001100000;
		sqrt_table[ 905] = 36'b111101001001110100000110100001011111;
		sqrt_table[ 906] = 36'b111101001100010000000000100001011110;
		sqrt_table[ 907] = 36'b111101001100110110111110100001011101;
		sqrt_table[ 908] = 36'b111101001111010011001100100001011100;
		sqrt_table[ 909] = 36'b111101010000100001010100100001011011;
		sqrt_table[ 910] = 36'b111101010001101111100010100001011011;
		sqrt_table[ 911] = 36'b111101010011100100111100100001011010;
		sqrt_table[ 912] = 36'b111101010101011010011100100001011001;
		sqrt_table[ 913] = 36'b111101010110101000110110100001011000;
		sqrt_table[ 914] = 36'b111101011000011110100010100001010111;
		sqrt_table[ 915] = 36'b111101011001101101000010100001010110;
		sqrt_table[ 916] = 36'b111101011011100010111000100001010101;
		sqrt_table[ 917] = 36'b111101011100110001100010100001010101;
		sqrt_table[ 918] = 36'b111101011110100111101000100001010100;
		sqrt_table[ 919] = 36'b111101100000011101110000100001010011;
		sqrt_table[ 920] = 36'b111101100001101100100110100001010010;
		sqrt_table[ 921] = 36'b111101100010111011011110100001010001;
		sqrt_table[ 922] = 36'b111101100100110001111100100001010000;
		sqrt_table[ 923] = 36'b111101100110101000011100100001001111;
		sqrt_table[ 924] = 36'b111101100111110111100010100001001111;
		sqrt_table[ 925] = 36'b111101101001101110010010100001001110;
		sqrt_table[ 926] = 36'b111101101010111101100010100001001101;
		sqrt_table[ 927] = 36'b111101101100001100110000100001001100;
		sqrt_table[ 928] = 36'b111101101110101011011100100001001011;
		sqrt_table[ 929] = 36'b111101101111010011001000100001001011;
		sqrt_table[ 930] = 36'b111101110001001010010100100001001010;
		sqrt_table[ 931] = 36'b111101110011000001100110100001001001;
		sqrt_table[ 932] = 36'b111101110100010001001100100001001000;
		sqrt_table[ 933] = 36'b111101110110001000101010100001000111;
		sqrt_table[ 934] = 36'b111101110111011000010110100001000110;
		sqrt_table[ 935] = 36'b111101111001001111111110100001000101;
		sqrt_table[ 936] = 36'b111101111010011111110100100001000101;
		sqrt_table[ 937] = 36'b111101111011101111101110100001000100;
		sqrt_table[ 938] = 36'b111101111101100111101100100001000011;
		sqrt_table[ 939] = 36'b111101111111011111101100100001000010;
		sqrt_table[ 940] = 36'b111110000000101111110000100001000001;
		sqrt_table[ 941] = 36'b111110000010101000000000100001000000;
		sqrt_table[ 942] = 36'b111110000011111000010000100001000000;
		sqrt_table[ 943] = 36'b111110000101001000100000100000111111;
		sqrt_table[ 944] = 36'b111110000111000000111110100000111110;
		sqrt_table[ 945] = 36'b111110001000010001010110100000111101;
		sqrt_table[ 946] = 36'b111110001010001010000100100000111100;
		sqrt_table[ 947] = 36'b111110001011011010100110100000111100;
		sqrt_table[ 948] = 36'b111110001101010011011110100000111011;
		sqrt_table[ 949] = 36'b111110001110100100001000100000111010;
		sqrt_table[ 950] = 36'b111110010000011101001100100000111001;
		sqrt_table[ 951] = 36'b111110010001101101111100100000111000;
		sqrt_table[ 952] = 36'b111110010011100111001010100000110111;
		sqrt_table[ 953] = 36'b111110010100111000000100100000110111;
		sqrt_table[ 954] = 36'b111110010110001001000010100000110110;
		sqrt_table[ 955] = 36'b111110011000000010100110100000110101;
		sqrt_table[ 956] = 36'b111110011001010011101010100000110100;
		sqrt_table[ 957] = 36'b111110011011001101011000100000110011;
		sqrt_table[ 958] = 36'b111110011100011110100110100000110011;
		sqrt_table[ 959] = 36'b111110011101101111111000100000110010;
		sqrt_table[ 960] = 36'b111110011111101001111000100000110001;
		sqrt_table[ 961] = 36'b111110100001100011111110100000110000;
		sqrt_table[ 962] = 36'b111110100010001100101100100000110000;
		sqrt_table[ 963] = 36'b111110100100101111101110100000101110;
		sqrt_table[ 964] = 36'b111110100101011000100010100000101110;
		sqrt_table[ 965] = 36'b111110100111010011000000100000101101;
		sqrt_table[ 966] = 36'b111110101000100100101100100000101100;
		sqrt_table[ 967] = 36'b111110101010011111010100100000101011;
		sqrt_table[ 968] = 36'b111110101011110001001010100000101011;
		sqrt_table[ 969] = 36'b111110101101101100000010100000101010;
		sqrt_table[ 970] = 36'b111110101110111110000000100000101001;
		sqrt_table[ 971] = 36'b111110110000010000000000100000101000;
		sqrt_table[ 972] = 36'b111110110010001011000110100000100111;
		sqrt_table[ 973] = 36'b111110110011011101010000100000100111;
		sqrt_table[ 974] = 36'b111110110101011000100110100000100110;
		sqrt_table[ 975] = 36'b111110110110101010111010100000100101;
		sqrt_table[ 976] = 36'b111110110111111101001100100000100100;
		sqrt_table[ 977] = 36'b111110111001001111100110100000100100;
		sqrt_table[ 978] = 36'b111110111011001011010010100000100011;
		sqrt_table[ 979] = 36'b111110111101000111000100100000100010;
		sqrt_table[ 980] = 36'b111110111110011001101010100000100001;
		sqrt_table[ 981] = 36'b111110111111101100010100100000100000;
		sqrt_table[ 982] = 36'b111111000000111111000000100000100000;
		sqrt_table[ 983] = 36'b111111000010111011001000100000011111;
		sqrt_table[ 984] = 36'b111111000100001101111110100000011110;
		sqrt_table[ 985] = 36'b111111000110001010010110100000011101;
		sqrt_table[ 986] = 36'b111111000110110011110100100000011101;
		sqrt_table[ 987] = 36'b111111001001011001110100100000011011;
		sqrt_table[ 988] = 36'b111111001010000011011010100000011011;
		sqrt_table[ 989] = 36'b111111001100000000001000100000011010;
		sqrt_table[ 990] = 36'b111111001101010011010100100000011001;
		sqrt_table[ 991] = 36'b111111001111010000001110100000011000;
		sqrt_table[ 992] = 36'b111111010000100011100100100000011000;
		sqrt_table[ 993] = 36'b111111010001110111000000100000010111;
		sqrt_table[ 994] = 36'b111111010011001010011010100000010110;
		sqrt_table[ 995] = 36'b111111010101000111101010100000010101;
		sqrt_table[ 996] = 36'b111111010110011011010000100000010101;
		sqrt_table[ 997] = 36'b111111011000011000110000100000010100;
		sqrt_table[ 998] = 36'b111111011001101100100000100000010011;
		sqrt_table[ 999] = 36'b111111011011000000001110100000010010;
		sqrt_table[1000] = 36'b111111011100010100000100100000010010;
		sqrt_table[1001] = 36'b111111011110010001111010100000010001;
		sqrt_table[1002] = 36'b111111011111100101111000100000010000;
		sqrt_table[1003] = 36'b111111100000111001111000100000001111;
		sqrt_table[1004] = 36'b111111100010111000000000100000001110;
		sqrt_table[1005] = 36'b111111100100001100001010100000001110;
		sqrt_table[1006] = 36'b111111100101100000011000100000001101;
		sqrt_table[1007] = 36'b111111100111011110110010100000001100;
		sqrt_table[1008] = 36'b111111101000110011000110100000001011;
		sqrt_table[1009] = 36'b111111101010000111100000100000001011;
		sqrt_table[1010] = 36'b111111101011011011111110100000001010;
		sqrt_table[1011] = 36'b111111101101011010110000100000001001;
		sqrt_table[1012] = 36'b111111101110101111010100100000001000;
		sqrt_table[1013] = 36'b111111110000000011111110100000001000;
		sqrt_table[1014] = 36'b111111110001011000101100100000000111;
		sqrt_table[1015] = 36'b111111110011010111110100100000000110;
		sqrt_table[1016] = 36'b111111110100101100101000100000000101;
		sqrt_table[1017] = 36'b111111110110101100000000100000000100;
		sqrt_table[1018] = 36'b111111110111010110100000100000000100;
		sqrt_table[1019] = 36'b111111111001010110000010100000000011;
		sqrt_table[1020] = 36'b111111111010101011000110100000000010;
		sqrt_table[1021] = 36'b111111111100101010110010100000000001;
		sqrt_table[1022] = 36'b111111111101010101011100100000000001;
		sqrt_table[1023] = 36'b111111111111010101010110100000000000;*/
	end
endmodule

`default_nettype wire