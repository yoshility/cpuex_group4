`default_nettype wire
module finv (
	input wire [31:0]  x,
  output wire [31:0] y,
  //output wire        ovf,
  input wire       clk,
  input wire       rstn
);
	wire      	sign = x[31];
	wire [ 7:0] exp_x = x[30:23];
	wire [22:0] frac_x = x[22:0];

	wire [ 9:0] addr = x[22:13];
	wire [12:0] dx = x[12:0];
	wire [35:0] dout;
	finv_table finv_table1(addr, dout, clk, rstn);

	wire [22:0] constant = dout[35:13];
	wire [12:0] gradient = dout[12:0];
	wire [25:0] dy_calc = gradient * dx;
	wire [23:0] frac_y = {constant,1'b0} - {10'b0, dy_calc[25:12]};

	wire [ 7:0] exp_y = 8'd253 - exp_x;

	assign y = {sign , exp_y, frac_y[22:0]};
endmodule

module fdiv (
	input  [31:0] x1,
	input  [31:0] x2,
	output [31:0] y,
	input 				clk,
	input					rstn
);
	wire [31:0] inv_x2;
	finv finv_in_fdiv(x2,inv_x2,clk,rstn);
	fmul fmul_in_fdiv(x1,inv_x2,y,clk,rstn);
endmodule

module finv_table (
	input		wire [ 9:0]	addr,
	output	reg  [35:0] dout,
	input 	wire 				clk,
	input 	wire 				rstn
);
	(*ram_style = "BLOCK"*) logic [35:0] finv_table [1023:0];
	always_comb begin
		dout = finv_table[addr];
	end
	initial begin
		finv_table[   0] = 36'b111111111111111111111111111111111000;
		finv_table[   1] = 36'b111111111100000000001111111111101000;
		finv_table[   2] = 36'b111111111000000000111111111111011000;
		finv_table[   3] = 36'b111111110100000010001111111111001000;
		finv_table[   4] = 36'b111111110000000011111101111110111000;
		finv_table[   5] = 36'b111111101100000110001101111110101000;
		finv_table[   6] = 36'b111111101000001000111011111110011000;
		finv_table[   7] = 36'b111111100100001100001001111110001001;
		finv_table[   8] = 36'b111111100000001111110101111101111001;
		finv_table[   9] = 36'b111111011100010100000011111101101010;
		finv_table[  10] = 36'b111111011000011000101111111101011010;
		finv_table[  11] = 36'b111111010100011101111001111101001011;
		finv_table[  12] = 36'b111111010000100011100011111100111011;
		finv_table[  13] = 36'b111111001100101001101101111100101100;
		finv_table[  14] = 36'b111111001000110000010011111100011100;
		finv_table[  15] = 36'b111111000100110111011011111100001101;
		finv_table[  16] = 36'b111111000000111110111111111011111110;
		finv_table[  17] = 36'b111110111101000111000011111011101111;
		finv_table[  18] = 36'b111110111001001111100101111011011111;
		finv_table[  19] = 36'b111110110101011000100101111011010000;
		finv_table[  20] = 36'b111110110001100010000011111011000001;
		finv_table[  21] = 36'b111110101101101100000001111010110010;
		finv_table[  22] = 36'b111110101001110110011011111010100011;
		finv_table[  23] = 36'b111110100110000001010101111010010100;
		finv_table[  24] = 36'b111110100010001100101011111010000101;
		finv_table[  25] = 36'b111110011110011000100001111001110110;
		finv_table[  26] = 36'b111110011010100100110011111001100111;
		finv_table[  27] = 36'b111110010110110001100011111001011001;
		finv_table[  28] = 36'b111110010010111110110001111001001010;
		finv_table[  29] = 36'b111110001111001100011011111000111011;
		finv_table[  30] = 36'b111110001011011010100101111000101100;
		finv_table[  31] = 36'b111110000111101001001011111000011110;
		finv_table[  32] = 36'b111110000011111000001101111000001111;
		finv_table[  33] = 36'b111110000000000111101111111000000001;
		finv_table[  34] = 36'b111101111100010111101011110111110010;
		finv_table[  35] = 36'b111101111000101000000111110111100100;
		finv_table[  36] = 36'b111101110100111000111101110111010101;
		finv_table[  37] = 36'b111101110001001010010011110111000111;
		finv_table[  38] = 36'b111101101101011100000011110110111001;
		finv_table[  39] = 36'b111101101001101110010001110110101010;
		finv_table[  40] = 36'b111101100110000000111101110110011100;
		finv_table[  41] = 36'b111101100010010100000011110110001110;
		finv_table[  42] = 36'b111101011110100111100111110110000000;
		finv_table[  43] = 36'b111101011010111011100101110101110001;
		finv_table[  44] = 36'b111101010111010000000011110101100011;
		finv_table[  45] = 36'b111101010011100100111011110101010101;
		finv_table[  46] = 36'b111101001111111010001111110101000111;
		finv_table[  47] = 36'b111101001100001111111111110100111001;
		finv_table[  48] = 36'b111101001000100110001011110100101011;
		finv_table[  49] = 36'b111101000100111100110011110100011101;
		finv_table[  50] = 36'b111101000001010011111001110100010000;
		finv_table[  51] = 36'b111100111101101011011001110100000010;
		finv_table[  52] = 36'b111100111010000011010011110011110100;
		finv_table[  53] = 36'b111100110110011011101011110011100110;
		finv_table[  54] = 36'b111100110010110100011101110011011000;
		finv_table[  55] = 36'b111100101111001101101011110011001011;
		finv_table[  56] = 36'b111100101011100111010101110010111101;
		finv_table[  57] = 36'b111100101000000001011001110010110000;
		finv_table[  58] = 36'b111100100100011011111001110010100010;
		finv_table[  59] = 36'b111100100000110110110011110010010100;
		finv_table[  60] = 36'b111100011101010010001011110010000111;
		finv_table[  61] = 36'b111100011001101101111011110001111010;
		finv_table[  62] = 36'b111100010110001010000111110001101100;
		finv_table[  63] = 36'b111100010010100110101101110001011111;
		finv_table[  64] = 36'b111100001111000011101111110001010001;
		finv_table[  65] = 36'b111100001011100001001011110001000100;
		finv_table[  66] = 36'b111100000111111111000011110000110111;
		finv_table[  67] = 36'b111100000100011101010101110000101010;
		finv_table[  68] = 36'b111100000000111011111111110000011100;
		finv_table[  69] = 36'b111011111101011011000101110000001111;
		finv_table[  70] = 36'b111011111001111010100111110000000010;
		finv_table[  71] = 36'b111011110110011010100001101111110101;
		finv_table[  72] = 36'b111011110010111010110101101111101000;
		finv_table[  73] = 36'b111011101111011011100101101111011011;
		finv_table[  74] = 36'b111011101011111100101101101111001110;
		finv_table[  75] = 36'b111011101000011110010001101111000001;
		finv_table[  76] = 36'b111011100101000000001101101110110100;
		finv_table[  77] = 36'b111011100001100010100011101110100111;
		finv_table[  78] = 36'b111011011110000101010101101110011010;
		finv_table[  79] = 36'b111011011010101000011111101110001110;
		finv_table[  80] = 36'b111011010111001100000011101110000001;
		finv_table[  81] = 36'b111011010011101111111111101101110100;
		finv_table[  82] = 36'b111011010000010100010101101101100111;
		finv_table[  83] = 36'b111011001100111001000111101101011011;
		finv_table[  84] = 36'b111011001001011110001111101101001110;
		finv_table[  85] = 36'b111011000110000011110011101101000010;
		finv_table[  86] = 36'b111011000010101001101111101100110101;
		finv_table[  87] = 36'b111010111111010000000011101100101000;
		finv_table[  88] = 36'b111010111011110110110001101100011100;
		finv_table[  89] = 36'b111010111000011101111001101100010000;
		finv_table[  90] = 36'b111010110101000101011001101100000011;
		finv_table[  91] = 36'b111010110001101101010001101011110111;
		finv_table[  92] = 36'b111010101110010101100011101011101010;
		finv_table[  93] = 36'b111010101010111110001101101011011110;
		finv_table[  94] = 36'b111010100111100111010001101011010010;
		finv_table[  95] = 36'b111010100100010000101011101011000101;
		finv_table[  96] = 36'b111010100000111010011111101010111001;
		finv_table[  97] = 36'b111010011101100100101101101010101101;
		finv_table[  98] = 36'b111010011010001111010001101010100001;
		finv_table[  99] = 36'b111010010110111010001111101010010101;
		finv_table[ 100] = 36'b111010010011100101100011101010001001;
				finv_table[ 101] = 36'b111010010000010001010001101001111101;
		finv_table[ 102] = 36'b111010001100111101010111101001110001;
		finv_table[ 103] = 36'b111010001001101001110111101001100101;
		finv_table[ 104] = 36'b111010000110010110101011101001011001;
		finv_table[ 105] = 36'b111010000011000011111001101001001101;
		finv_table[ 106] = 36'b111001111111110001011111101001000001;
		finv_table[ 107] = 36'b111001111100011111011101101000110101;
		finv_table[ 108] = 36'b111001111001001101110001101000101001;
		finv_table[ 109] = 36'b111001110101111100011111101000011101;
		finv_table[ 110] = 36'b111001110010101011100011101000010001;
		finv_table[ 111] = 36'b111001101111011011000001101000000110;
		finv_table[ 112] = 36'b111001101100001010110011100111111010;
		finv_table[ 113] = 36'b111001101000111010111111100111101110;
		finv_table[ 114] = 36'b111001100101101011100001100111100011;
		finv_table[ 115] = 36'b111001100010011100011011100111010111;
		finv_table[ 116] = 36'b111001011111001101101011100111001011;
		finv_table[ 117] = 36'b111001011011111111010101100111000000;
		finv_table[ 118] = 36'b111001011000110001010011100110110100;
		finv_table[ 119] = 36'b111001010101100011101011100110101001;
		finv_table[ 120] = 36'b111001010010010110010111100110011101;
		finv_table[ 121] = 36'b111001001111001001011011100110010010;
		finv_table[ 122] = 36'b111001001011111100110111100110000110;
		finv_table[ 123] = 36'b111001001000110000101001100101111011;
		finv_table[ 124] = 36'b111001000101100100110011100101110000;
		finv_table[ 125] = 36'b111001000010011001010001100101100100;
		finv_table[ 126] = 36'b111000111111001110000111100101011001;
		finv_table[ 127] = 36'b111000111100000011010101100101001110;
		finv_table[ 128] = 36'b111000111000111000110111100101000011;
		finv_table[ 129] = 36'b111000110101101110110001100100110111;
		finv_table[ 130] = 36'b111000110010100101000001100100101100;
		finv_table[ 131] = 36'b111000101111011011101001100100100001;
		finv_table[ 132] = 36'b111000101100010010100101100100010110;
		finv_table[ 133] = 36'b111000101001001001111001100100001011;
		finv_table[ 134] = 36'b111000100110000001100011100100000000;
		finv_table[ 135] = 36'b111000100010111001100011100011110101;
		finv_table[ 136] = 36'b111000011111110001110111100011101010;
		finv_table[ 137] = 36'b111000011100101010100011100011011111;
		finv_table[ 138] = 36'b111000011001100011100101100011010100;
		finv_table[ 139] = 36'b111000010110011100111011100011001001;
		finv_table[ 140] = 36'b111000010011010110101001100010111110;
		finv_table[ 141] = 36'b111000010000010000101011100010110011;
		finv_table[ 142] = 36'b111000001101001011000101100010101000;
		finv_table[ 143] = 36'b111000001010000101110011100010011101;
		finv_table[ 144] = 36'b111000000111000000110111100010010011;
		finv_table[ 145] = 36'b111000000011111100010001100010001000;
		finv_table[ 146] = 36'b111000000000110111111111100001111101;
		finv_table[ 147] = 36'b110111111101110100000101100001110011;
		finv_table[ 148] = 36'b110111111010110000011111100001101000;
		finv_table[ 149] = 36'b110111110111101101001101100001011101;
		finv_table[ 150] = 36'b110111110100101010010011100001010011;
		finv_table[ 151] = 36'b110111110001100111101101100001001000;
		finv_table[ 152] = 36'b110111101110100101011011100000111101;
		finv_table[ 153] = 36'b110111101011100011011111100000110011;
		finv_table[ 154] = 36'b110111101000100001111001100000101000;
		finv_table[ 155] = 36'b110111100101100000100111100000011110;
		finv_table[ 156] = 36'b110111100010011111101011100000010011;
		finv_table[ 157] = 36'b110111011111011111000011100000001001;
		finv_table[ 158] = 36'b110111011100011110101111011111111111;
		finv_table[ 159] = 36'b110111011001011110110001011111110100;
		finv_table[ 160] = 36'b110111010110011111001001011111101010;
		finv_table[ 161] = 36'b110111010011011111110011011111100000;
		finv_table[ 162] = 36'b110111010000100000110011011111010101;
		finv_table[ 163] = 36'b110111001101100010000111011111001011;
		finv_table[ 164] = 36'b110111001010100011110001011111000001;
		finv_table[ 165] = 36'b110111000111100101101101011110110111;
		finv_table[ 166] = 36'b110111000100100111111111011110101100;
		finv_table[ 167] = 36'b110111000001101010100111011110100010;
		finv_table[ 168] = 36'b110110111110101101100001011110011000;
		finv_table[ 169] = 36'b110110111011110000110001011110001110;
		finv_table[ 170] = 36'b110110111000110100010011011110000100;
		finv_table[ 171] = 36'b110110110101111000001011011101111010;
		finv_table[ 172] = 36'b110110110010111100010111011101110000;
		finv_table[ 173] = 36'b110110110000000000110111011101100110;
		finv_table[ 174] = 36'b110110101101000101101001011101011100;
		finv_table[ 175] = 36'b110110101010001010110001011101010010;
		finv_table[ 176] = 36'b110110100111010000001101011101001000;
		finv_table[ 177] = 36'b110110100100010101111101011100111110;
		finv_table[ 178] = 36'b110110100001011011111111011100110100;
		finv_table[ 179] = 36'b110110011110100010010111011100101010;
		finv_table[ 180] = 36'b110110011011101001000001011100100000;
		finv_table[ 181] = 36'b110110011000101111111111011100010110;
		finv_table[ 182] = 36'b110110010101110111010001011100001101;
		finv_table[ 183] = 36'b110110010010111110111001011100000011;
		finv_table[ 184] = 36'b110110010000000110110001011011111001;
		finv_table[ 185] = 36'b110110001101001110111101011011101111;
		finv_table[ 186] = 36'b110110001010010111011111011011100110;
		finv_table[ 187] = 36'b110110000111100000010011011011011100;
		finv_table[ 188] = 36'b110110000100101001011001011011010010;
		finv_table[ 189] = 36'b110110000001110010110011011011001001;
		finv_table[ 190] = 36'b110101111110111100100001011010111111;
		finv_table[ 191] = 36'b110101111100000110100001011010110110;
		finv_table[ 192] = 36'b110101111001010000110101011010101100;
		finv_table[ 193] = 36'b110101110110011011011011011010100010;
		finv_table[ 194] = 36'b110101110011100110010111011010011001;
		finv_table[ 195] = 36'b110101110000110001100011011010001111;
		finv_table[ 196] = 36'b110101101101111101000011011010000110;
		finv_table[ 197] = 36'b110101101011001000110101011001111101;
		finv_table[ 198] = 36'b110101101000010100111101011001110011;
		finv_table[ 199] = 36'b110101100101100001010101011001101010;
		finv_table[ 200] = 36'b110101100010101110000001011001100000;
		finv_table[ 201] = 36'b110101011111111010111111011001010111;
		finv_table[ 202] = 36'b110101011101001000001111011001001110;
		finv_table[ 203] = 36'b110101011010010101110011011001000100;
		finv_table[ 204] = 36'b110101010111100011101001011000111011;
		finv_table[ 205] = 36'b110101010100110001110001011000110010;
		finv_table[ 206] = 36'b110101010010000000001101011000101001;
		finv_table[ 207] = 36'b110101001111001110111011011000011111;
		finv_table[ 208] = 36'b110101001100011101111011011000010110;
		finv_table[ 209] = 36'b110101001001101101001101011000001101;
		finv_table[ 210] = 36'b110101000110111100110001011000000100;
		finv_table[ 211] = 36'b110101000100001100101001010111111011;
		finv_table[ 212] = 36'b110101000001011100110011010111110010;
		finv_table[ 213] = 36'b110100111110101101001101010111101001;
		finv_table[ 214] = 36'b110100111011111101111011010111100000;
		finv_table[ 215] = 36'b110100111001001110111011010111010111;
		finv_table[ 216] = 36'b110100110110100000001101010111001110;
		finv_table[ 217] = 36'b110100110011110001110001010111000101;
		finv_table[ 218] = 36'b110100110001000011100111010110111100;
		finv_table[ 219] = 36'b110100101110010101101111010110110011;
		finv_table[ 220] = 36'b110100101011101000000111010110101010;
		finv_table[ 221] = 36'b110100101000111010110011010110100001;
		finv_table[ 222] = 36'b110100100110001101110001010110011000;
		finv_table[ 223] = 36'b110100100011100000111111010110001111;
		finv_table[ 224] = 36'b110100100000110100100001010110000110;
		finv_table[ 225] = 36'b110100011110001000010011010101111101;
		finv_table[ 226] = 36'b110100011011011100010111010101110101;
		finv_table[ 227] = 36'b110100011000110000101101010101101100;
		finv_table[ 228] = 36'b110100010110000101010011010101100011;
		finv_table[ 229] = 36'b110100010011011010001101010101011010;
		finv_table[ 230] = 36'b110100010000101111010111010101010010;
		finv_table[ 231] = 36'b110100001110000100110011010101001001;
		finv_table[ 232] = 36'b110100001011011010011111010101000000;
		finv_table[ 233] = 36'b110100001000110000011101010100111000;
		finv_table[ 234] = 36'b110100000110000110101101010100101111;
		finv_table[ 235] = 36'b110100000011011101001111010100100110;
		finv_table[ 236] = 36'b110100000000110100000001010100011110;
		finv_table[ 237] = 36'b110011111110001011000011010100010101;
		finv_table[ 238] = 36'b110011111011100010011001010100001101;
		finv_table[ 239] = 36'b110011111000111001111101010100000100;
		finv_table[ 240] = 36'b110011110110010001110101010011111100;
		finv_table[ 241] = 36'b110011110011101001111011010011110011;
		finv_table[ 242] = 36'b110011110001000010010101010011101011;
		finv_table[ 243] = 36'b110011101110011010111101010011100010;
		finv_table[ 244] = 36'b110011101011110011111001010011011010;
		finv_table[ 245] = 36'b110011101001001101000011010011010001;
		finv_table[ 246] = 36'b110011100110100110011111010011001001;
		finv_table[ 247] = 36'b110011100100000000001101010011000001;
		finv_table[ 248] = 36'b110011100001011010001001010010111000;
		finv_table[ 249] = 36'b110011011110110100011001010010110000;
		finv_table[ 250] = 36'b110011011100001110110111010010101000;
		finv_table[ 251] = 36'b110011011001101001100111010010011111;
		finv_table[ 252] = 36'b110011010111000100100111010010010111;
		finv_table[ 253] = 36'b110011010100011111110111010010001111;
		finv_table[ 254] = 36'b110011010001111011011001010010000111;
		finv_table[ 255] = 36'b110011001111010111001011010001111110;
		finv_table[ 256] = 36'b110011001100110011001101010001110110;
		finv_table[ 257] = 36'b110011001010001111011111010001101110;
		finv_table[ 258] = 36'b110011000111101100000001010001100110;
		finv_table[ 259] = 36'b110011000101001000110101010001011110;
		finv_table[ 260] = 36'b110011000010100101110111010001010110;
		finv_table[ 261] = 36'b110011000000000011001011010001001110;
		finv_table[ 262] = 36'b110010111101100000101111010001000110;
		finv_table[ 263] = 36'b110010111010111110100011010000111101;
		finv_table[ 264] = 36'b110010111000011100100111010000110101;
		finv_table[ 265] = 36'b110010110101111010111011010000101101;
		finv_table[ 266] = 36'b110010110011011001011111010000100101;
		finv_table[ 267] = 36'b110010110000111000010011010000011101;
		finv_table[ 268] = 36'b110010101110010111010111010000010101;
		finv_table[ 269] = 36'b110010101011110110101011010000001110;
		finv_table[ 270] = 36'b110010101001010110001111010000000110;
		finv_table[ 271] = 36'b110010100110110110000011001111111110;
		finv_table[ 272] = 36'b110010100100010110001001001111110110;
		finv_table[ 273] = 36'b110010100001110110011011001111101110;
		finv_table[ 274] = 36'b110010011111010110111111001111100110;
		finv_table[ 275] = 36'b110010011100110111110001001111011110;
		finv_table[ 276] = 36'b110010011010011000110011001111010110;
		finv_table[ 277] = 36'b110010010111111010000101001111001111;
		finv_table[ 278] = 36'b110010010101011011101001001111000111;
		finv_table[ 279] = 36'b110010010010111101011001001110111111;
		finv_table[ 280] = 36'b110010010000011111011001001110110111;
		finv_table[ 281] = 36'b110010001110000001101011001110110000;
		finv_table[ 282] = 36'b110010001011100100001011001110101000;
		finv_table[ 283] = 36'b110010001001000110111001001110100000;
		finv_table[ 284] = 36'b110010000110101001111001001110011000;
		finv_table[ 285] = 36'b110010000100001101000111001110010001;
		finv_table[ 286] = 36'b110010000001110000100011001110001001;
		finv_table[ 287] = 36'b110001111111010100010001001110000010;
		finv_table[ 288] = 36'b110001111100111000001011001101111010;
		finv_table[ 289] = 36'b110001111010011100010111001101110010;
		finv_table[ 290] = 36'b110001111000000000110011001101101011;
		finv_table[ 291] = 36'b110001110101100101011011001101100011;
		finv_table[ 292] = 36'b110001110011001010010101001101011100;
		finv_table[ 293] = 36'b110001110000101111011011001101010100;
		finv_table[ 294] = 36'b110001101110010100110001001101001101;
		finv_table[ 295] = 36'b110001101011111010010111001101000101;
		finv_table[ 296] = 36'b110001101001100000001011001100111110;
		finv_table[ 297] = 36'b110001100111000110001111001100110110;
		finv_table[ 298] = 36'b110001100100101100100001001100101111;
		finv_table[ 299] = 36'b110001100010010011000011001100100111;
		finv_table[ 300] = 36'b110001011111111001110101001100100000;
		finv_table[ 301] = 36'b110001011101100000110011001100011001;
		finv_table[ 302] = 36'b110001011011001000000001001100010001;
		finv_table[ 303] = 36'b110001011000101111011101001100001010;
		finv_table[ 304] = 36'b110001010110010111000111001100000011;
		finv_table[ 305] = 36'b110001010011111111000011001011111011;
		finv_table[ 306] = 36'b110001010001100111001011001011110100;
		finv_table[ 307] = 36'b110001001111001111100001001011101101;
		finv_table[ 308] = 36'b110001001100111000000111001011100101;
		finv_table[ 309] = 36'b110001001010100000111011001011011110;
		finv_table[ 310] = 36'b110001001000001001111111001011010111;
		finv_table[ 311] = 36'b110001000101110011001111001011010000;
		finv_table[ 312] = 36'b110001000011011100101111001011001000;
		finv_table[ 313] = 36'b110001000001000110011101001011000001;
		finv_table[ 314] = 36'b110000111110110000011011001010111010;
		finv_table[ 315] = 36'b110000111100011010100101001010110011;
		finv_table[ 316] = 36'b110000111010000100111111001010101100;
		finv_table[ 317] = 36'b110000110111101111100101001010100101;
		finv_table[ 318] = 36'b110000110101011010011011001010011110;
		finv_table[ 319] = 36'b110000110011000101011111001010010110;
		finv_table[ 320] = 36'b110000110000110000110001001010001111;
		finv_table[ 321] = 36'b110000101110011100010001001010001000;
		finv_table[ 322] = 36'b110000101100000111111111001010000001;
		finv_table[ 323] = 36'b110000101001110011111011001001111010;
		finv_table[ 324] = 36'b110000100111100000000101001001110011;
		finv_table[ 325] = 36'b110000100101001100011111001001101100;
		finv_table[ 326] = 36'b110000100010111001000101001001100101;
		finv_table[ 327] = 36'b110000100000100101111001001001011110;
		finv_table[ 328] = 36'b110000011110010010111011001001010111;
		finv_table[ 329] = 36'b110000011100000000001011001001010000;
		finv_table[ 330] = 36'b110000011001101101101011001001001010;
		finv_table[ 331] = 36'b110000010111011011010101001001000011;
		finv_table[ 332] = 36'b110000010101001001001111001000111100;
		finv_table[ 333] = 36'b110000010010110111011001001000110101;
		finv_table[ 334] = 36'b110000010000100101101101001000101110;
		finv_table[ 335] = 36'b110000001110010100010001001000100111;
		finv_table[ 336] = 36'b110000001100000011000001001000100000;
		finv_table[ 337] = 36'b110000001001110001111111001000011001;
		finv_table[ 338] = 36'b110000000111100001001011001000010011;
		finv_table[ 339] = 36'b110000000101010000100101001000001100;
		finv_table[ 340] = 36'b110000000011000000001101001000000101;
		finv_table[ 341] = 36'b110000000000110000000001000111111110;
		finv_table[ 342] = 36'b101111111110100000000011000111111000;
		finv_table[ 343] = 36'b101111111100010000010011000111110001;
		finv_table[ 344] = 36'b101111111010000000101111000111101010;
		finv_table[ 345] = 36'b101111110111110001011011000111100100;
		finv_table[ 346] = 36'b101111110101100010010001000111011101;
		finv_table[ 347] = 36'b101111110011010011010111000111010110;
		finv_table[ 348] = 36'b101111110001000100101011000111010000;
		finv_table[ 349] = 36'b101111101110110110001011000111001001;
		finv_table[ 350] = 36'b101111101100100111110111000111000010;
		finv_table[ 351] = 36'b101111101010011001110011000110111100;
		finv_table[ 352] = 36'b101111101000001011111011000110110101;
		finv_table[ 353] = 36'b101111100101111110001111000110101110;
		finv_table[ 354] = 36'b101111100011110000110001000110101000;
		finv_table[ 355] = 36'b101111100001100011100001000110100001;
		finv_table[ 356] = 36'b101111011111010110011101000110011011;
		finv_table[ 357] = 36'b101111011101001001100101000110010100;
		finv_table[ 358] = 36'b101111011010111100111011000110001110;
		finv_table[ 359] = 36'b101111011000110000011111000110000111;
		finv_table[ 360] = 36'b101111010110100100001111000110000001;
		finv_table[ 361] = 36'b101111010100011000001101000101111010;
		finv_table[ 362] = 36'b101111010010001100011001000101110100;
		finv_table[ 363] = 36'b101111010000000000101111000101101101;
		finv_table[ 364] = 36'b101111001101110101010011000101100111;
		finv_table[ 365] = 36'b101111001011101010000011000101100001;
		finv_table[ 366] = 36'b101111001001011111000011000101011010;
		finv_table[ 367] = 36'b101111000111010100001101000101010100;
		finv_table[ 368] = 36'b101111000101001001100011000101001101;
		finv_table[ 369] = 36'b101111000010111111001001000101000111;
		finv_table[ 370] = 36'b101111000000110100111001000101000001;
		finv_table[ 371] = 36'b101110111110101010110111000100111010;
		finv_table[ 372] = 36'b101110111100100001000001000100110100;
		finv_table[ 373] = 36'b101110111010010111010111000100101110;
		finv_table[ 374] = 36'b101110111000001101111011000100101000;
		finv_table[ 375] = 36'b101110110110000100101011000100100001;
		finv_table[ 376] = 36'b101110110011111011100111000100011011;
		finv_table[ 377] = 36'b101110110001110010101111000100010101;
		finv_table[ 378] = 36'b101110101111101010000101000100001111;
		finv_table[ 379] = 36'b101110101101100001100111000100001000;
		finv_table[ 380] = 36'b101110101011011001010111000100000010;
		finv_table[ 381] = 36'b101110101001010001010001000011111100;
		finv_table[ 382] = 36'b101110100111001001010111000011110110;
		finv_table[ 383] = 36'b101110100101000001101011000011110000;
		finv_table[ 384] = 36'b101110100010111010001011000011101001;
		finv_table[ 385] = 36'b101110100000110010111001000011100011;
		finv_table[ 386] = 36'b101110011110101011110001000011011101;
		finv_table[ 387] = 36'b101110011100100100110101000011010111;
		finv_table[ 388] = 36'b101110011010011110000111000011010001;
		finv_table[ 389] = 36'b101110011000010111100011000011001011;
		finv_table[ 390] = 36'b101110010110010001001101000011000101;
		finv_table[ 391] = 36'b101110010100001011000001000010111111;
		finv_table[ 392] = 36'b101110010010000101000011000010111001;
		finv_table[ 393] = 36'b101110001111111111010001000010110011;
		finv_table[ 394] = 36'b101110001101111001101101000010101101;
		finv_table[ 395] = 36'b101110001011110100010001000010100111;
		finv_table[ 396] = 36'b101110001001101111000011000010100001;
		finv_table[ 397] = 36'b101110000111101010000001000010011011;
		finv_table[ 398] = 36'b101110000101100101001011000010010101;
		finv_table[ 399] = 36'b101110000011100000100001000010001111;
		finv_table[ 400] = 36'b101110000001011100000011000010001001;
				finv_table[ 401] = 36'b101101111111010111110001000010000011;
		finv_table[ 402] = 36'b101101111101010011101011000001111101;
		finv_table[ 403] = 36'b101101111011001111101111000001110111;
		finv_table[ 404] = 36'b101101111001001100000001000001110001;
		finv_table[ 405] = 36'b101101110111001000011111000001101011;
		finv_table[ 406] = 36'b101101110101000101000111000001100101;
		finv_table[ 407] = 36'b101101110011000001111011000001011111;
		finv_table[ 408] = 36'b101101110000111110111011000001011010;
		finv_table[ 409] = 36'b101101101110111100000111000001010100;
		finv_table[ 410] = 36'b101101101100111001011111000001001110;
		finv_table[ 411] = 36'b101101101010110111000011000001001000;
		finv_table[ 412] = 36'b101101101000110100110001000001000010;
		finv_table[ 413] = 36'b101101100110110010101011000000111100;
		finv_table[ 414] = 36'b101101100100110000110001000000110111;
		finv_table[ 415] = 36'b101101100010101111000101000000110001;
		finv_table[ 416] = 36'b101101100000101101100001000000101011;
		finv_table[ 417] = 36'b101101011110101100001001000000100101;
		finv_table[ 418] = 36'b101101011100101010111111000000100000;
		finv_table[ 419] = 36'b101101011010101001111101000000011010;
		finv_table[ 420] = 36'b101101011000101001001001000000010100;
		finv_table[ 421] = 36'b101101010110101000011111000000001111;
		finv_table[ 422] = 36'b101101010100101000000001000000001001;
		finv_table[ 423] = 36'b101101010010100111101111000000000011;
		finv_table[ 424] = 36'b101101010000100111100110111111111110;
		finv_table[ 425] = 36'b101101001110100111101010111111111000;
		finv_table[ 426] = 36'b101101001100100111111000111111110010;
		finv_table[ 427] = 36'b101101001010101000010010111111101101;
		finv_table[ 428] = 36'b101101001000101000111010111111100111;
		finv_table[ 429] = 36'b101101000110101001101010111111100001;
		finv_table[ 430] = 36'b101101000100101010100110111111011100;
		finv_table[ 431] = 36'b101101000010101011101110111111010110;
		finv_table[ 432] = 36'b101101000000101101000000111111010001;
		finv_table[ 433] = 36'b101100111110101110011110111111001011;
		finv_table[ 434] = 36'b101100111100110000000110111111000110;
		finv_table[ 435] = 36'b101100111010110001111010111111000000;
		finv_table[ 436] = 36'b101100111000110011111000111110111011;
		finv_table[ 437] = 36'b101100110110110110000100111110110101;
		finv_table[ 438] = 36'b101100110100111000011000111110110000;
		finv_table[ 439] = 36'b101100110010111010111000111110101010;
		finv_table[ 440] = 36'b101100110000111101100010111110100101;
		finv_table[ 441] = 36'b101100101111000000011000111110011111;
		finv_table[ 442] = 36'b101100101101000011011000111110011010;
		finv_table[ 443] = 36'b101100101011000110100100111110010100;
		finv_table[ 444] = 36'b101100101001001001111010111110001111;
		finv_table[ 445] = 36'b101100100111001101011100111110001001;
		finv_table[ 446] = 36'b101100100101010001001010111110000100;
		finv_table[ 447] = 36'b101100100011010101000000111101111111;
		finv_table[ 448] = 36'b101100100001011001000010111101111001;
		finv_table[ 449] = 36'b101100011111011101001110111101110100;
		finv_table[ 450] = 36'b101100011101100001100110111101101110;
		finv_table[ 451] = 36'b101100011011100110001000111101101001;
		finv_table[ 452] = 36'b101100011001101010110110111101100100;
		finv_table[ 453] = 36'b101100010111101111101100111101011110;
		finv_table[ 454] = 36'b101100010101110100101110111101011001;
		finv_table[ 455] = 36'b101100010011111001111100111101010100;
		finv_table[ 456] = 36'b101100010001111111010010111101001110;
		finv_table[ 457] = 36'b101100010000000100110110111101001001;
		finv_table[ 458] = 36'b101100001110001010100010111101000100;
		finv_table[ 459] = 36'b101100001100010000011010111100111111;
		finv_table[ 460] = 36'b101100001010010110011010111100111001;
		finv_table[ 461] = 36'b101100001000011100100110111100110100;
		finv_table[ 462] = 36'b101100000110100010111110111100101111;
		finv_table[ 463] = 36'b101100000100101001011110111100101010;
		finv_table[ 464] = 36'b101100000010110000001010111100100100;
		finv_table[ 465] = 36'b101100000000110111000000111100011111;
		finv_table[ 466] = 36'b101011111110111110000000111100011010;
		finv_table[ 467] = 36'b101011111101000101001010111100010101;
		finv_table[ 468] = 36'b101011111011001100100010111100010000;
		finv_table[ 469] = 36'b101011111001010100000000111100001011;
		finv_table[ 470] = 36'b101011110111011011101010111100000101;
		finv_table[ 471] = 36'b101011110101100011011110111100000000;
		finv_table[ 472] = 36'b101011110011101011011110111011111011;
		finv_table[ 473] = 36'b101011110001110011100110111011110110;
		finv_table[ 474] = 36'b101011101111111011111010111011110001;
		finv_table[ 475] = 36'b101011101110000100010110111011101100;
		finv_table[ 476] = 36'b101011101100001100111100111011100111;
		finv_table[ 477] = 36'b101011101010010101110000111011100010;
		finv_table[ 478] = 36'b101011101000011110101010111011011101;
		finv_table[ 479] = 36'b101011100110100111110000111011010111;
		finv_table[ 480] = 36'b101011100100110001000000111011010010;
		finv_table[ 481] = 36'b101011100010111010011010111011001101;
		finv_table[ 482] = 36'b101011100001000011111110111011001000;
		finv_table[ 483] = 36'b101011011111001101101110111011000011;
		finv_table[ 484] = 36'b101011011101010111100110111010111110;
		finv_table[ 485] = 36'b101011011011100001101000111010111001;
		finv_table[ 486] = 36'b101011011001101011110100111010110100;
		finv_table[ 487] = 36'b101011010111110110001010111010101111;
		finv_table[ 488] = 36'b101011010110000000101010111010101010;
		finv_table[ 489] = 36'b101011010100001011010100111010100101;
		finv_table[ 490] = 36'b101011010010010110001000111010100000;
		finv_table[ 491] = 36'b101011010000100001000110111010011100;
		finv_table[ 492] = 36'b101011001110101100010000111010010111;
		finv_table[ 493] = 36'b101011001100110111100000111010010010;
		finv_table[ 494] = 36'b101011001011000010111100111010001101;
		finv_table[ 495] = 36'b101011001001001110100010111010001000;
		finv_table[ 496] = 36'b101011000111011010010010111010000011;
		finv_table[ 497] = 36'b101011000101100110001010111001111110;
		finv_table[ 498] = 36'b101011000011110010001100111001111001;
		finv_table[ 499] = 36'b101011000001111110011000111001110100;
		finv_table[ 500] = 36'b101011000000001010110000111001110000;
		finv_table[ 501] = 36'b101010111110010111001110111001101011;
		finv_table[ 502] = 36'b101010111100100011111010111001100110;
		finv_table[ 503] = 36'b101010111010110000101100111001100001;
		finv_table[ 504] = 36'b101010111000111101101000111001011100;
		finv_table[ 505] = 36'b101010110111001010110000111001010111;
		finv_table[ 506] = 36'b101010110101011000000000111001010011;
		finv_table[ 507] = 36'b101010110011100101011010111001001110;
		finv_table[ 508] = 36'b101010110001110010111110111001001001;
		finv_table[ 509] = 36'b101010110000000000101010111001000100;
		finv_table[ 510] = 36'b101010101110001110100000111001000000;
		finv_table[ 511] = 36'b101010101100011100100000111000111011;
		finv_table[ 512] = 36'b101010101010101010101010111000110110;
		finv_table[ 513] = 36'b101010101000111000111110111000110001;
		finv_table[ 514] = 36'b101010100111000111011000111000101101;
		finv_table[ 515] = 36'b101010100101010110000000111000101000;
		finv_table[ 516] = 36'b101010100011100100101110111000100011;
		finv_table[ 517] = 36'b101010100001110011100110111000011110;
		finv_table[ 518] = 36'b101010100000000010101010111000011010;
		finv_table[ 519] = 36'b101010011110010001110110111000010101;
		finv_table[ 520] = 36'b101010011100100001001000111000010000;
		finv_table[ 521] = 36'b101010011010110000101000111000001100;
		finv_table[ 522] = 36'b101010011001000000010000111000000111;
		finv_table[ 523] = 36'b101010010111010000000000111000000010;
		finv_table[ 524] = 36'b101010010101011111111010110111111110;
		finv_table[ 525] = 36'b101010010011101111111110110111111001;
		finv_table[ 526] = 36'b101010010010000000001010110111110101;
		finv_table[ 527] = 36'b101010010000010000100000110111110000;
		finv_table[ 528] = 36'b101010001110100000111110110111101011;
		finv_table[ 529] = 36'b101010001100110001101000110111100111;
		finv_table[ 530] = 36'b101010001011000010011000110111100010;
		finv_table[ 531] = 36'b101010001001010011010010110111011110;
		finv_table[ 532] = 36'b101010000111100100010110110111011001;
		finv_table[ 533] = 36'b101010000101110101100010110111010101;
		finv_table[ 534] = 36'b101010000100000110111010110111010000;
		finv_table[ 535] = 36'b101010000010011000011000110111001011;
		finv_table[ 536] = 36'b101010000000101010000000110111000111;
		finv_table[ 537] = 36'b101001111110111011110000110111000010;
		finv_table[ 538] = 36'b101001111101001101101100110110111110;
		finv_table[ 539] = 36'b101001111011011111101110110110111001;
		finv_table[ 540] = 36'b101001111001110001111010110110110101;
		finv_table[ 541] = 36'b101001111000000100001110110110110000;
		finv_table[ 542] = 36'b101001110110010110101110110110101100;
		finv_table[ 543] = 36'b101001110100101001010100110110101000;
		finv_table[ 544] = 36'b101001110010111100000100110110100011;
		finv_table[ 545] = 36'b101001110001001110111100110110011111;
		finv_table[ 546] = 36'b101001101111100001111110110110011010;
		finv_table[ 547] = 36'b101001101101110101001010110110010110;
		finv_table[ 548] = 36'b101001101100001000011110110110010001;
		finv_table[ 549] = 36'b101001101010011011111010110110001101;
		finv_table[ 550] = 36'b101001101000101111011110110110001001;
		finv_table[ 551] = 36'b101001100111000011001100110110000100;
		finv_table[ 552] = 36'b101001100101010111000100110110000000;
		finv_table[ 553] = 36'b101001100011101011000100110101111011;
		finv_table[ 554] = 36'b101001100001111111001100110101110111;
		finv_table[ 555] = 36'b101001100000010011011100110101110011;
		finv_table[ 556] = 36'b101001011110100111110110110101101110;
		finv_table[ 557] = 36'b101001011100111100011000110101101010;
		finv_table[ 558] = 36'b101001011011010001000100110101100110;
		finv_table[ 559] = 36'b101001011001100101111000110101100001;
		finv_table[ 560] = 36'b101001010111111010110100110101011101;
		finv_table[ 561] = 36'b101001010110001111111000110101011001;
		finv_table[ 562] = 36'b101001010100100101000110110101010100;
		finv_table[ 563] = 36'b101001010010111010011110110101010000;
		finv_table[ 564] = 36'b101001010001001111111100110101001100;
		finv_table[ 565] = 36'b101001001111100101100100110101000111;
		finv_table[ 566] = 36'b101001001101111011010100110101000011;
		finv_table[ 567] = 36'b101001001100010001001110110100111111;
		finv_table[ 568] = 36'b101001001010100111001110110100111011;
		finv_table[ 569] = 36'b101001001000111101011000110100110110;
		finv_table[ 570] = 36'b101001000111010011101010110100110010;
		finv_table[ 571] = 36'b101001000101101010000110110100101110;
		finv_table[ 572] = 36'b101001000100000000101000110100101010;
		finv_table[ 573] = 36'b101001000010010111010100110100100101;
		finv_table[ 574] = 36'b101001000000101110001000110100100001;
		finv_table[ 575] = 36'b101000111111000101000110110100011101;
		finv_table[ 576] = 36'b101000111101011100001000110100011001;
		finv_table[ 577] = 36'b101000111011110011011000110100010101;
		finv_table[ 578] = 36'b101000111010001010101100110100010000;
		finv_table[ 579] = 36'b101000111000100010001010110100001100;
		finv_table[ 580] = 36'b101000110110111001110000110100001000;
		finv_table[ 581] = 36'b101000110101010001100000110100000100;
		finv_table[ 582] = 36'b101000110011101001010110110100000000;
		finv_table[ 583] = 36'b101000110010000001010110110011111100;
		finv_table[ 584] = 36'b101000110000011001011110110011111000;
		finv_table[ 585] = 36'b101000101110110001101110110011110011;
		finv_table[ 586] = 36'b101000101101001010000110110011101111;
		finv_table[ 587] = 36'b101000101011100010100110110011101011;
		finv_table[ 588] = 36'b101000101001111011001110110011100111;
		finv_table[ 589] = 36'b101000101000010100000000110011100011;
		finv_table[ 590] = 36'b101000100110101100111000110011011111;
		finv_table[ 591] = 36'b101000100101000101111010110011011011;
		finv_table[ 592] = 36'b101000100011011111000010110011010111;
		finv_table[ 593] = 36'b101000100001111000010100110011010011;
		finv_table[ 594] = 36'b101000100000010001101100110011001111;
		finv_table[ 595] = 36'b101000011110101011001110110011001011;
		finv_table[ 596] = 36'b101000011101000100111010110011000111;
		finv_table[ 597] = 36'b101000011011011110101010110011000011;
		finv_table[ 598] = 36'b101000011001111000100100110010111111;
		finv_table[ 599] = 36'b101000011000010010100110110010111011;
		finv_table[ 600] = 36'b101000010110101100110000110010110110;
		finv_table[ 601] = 36'b101000010101000111000010110010110010;
		finv_table[ 602] = 36'b101000010011100001011100110010101110;
		finv_table[ 603] = 36'b101000010001111011111110110010101011;
		finv_table[ 604] = 36'b101000010000010110101000110010100111;
		finv_table[ 605] = 36'b101000001110110001011010110010100011;
		finv_table[ 606] = 36'b101000001101001100010100110010011111;
		finv_table[ 607] = 36'b101000001011100111010110110010011011;
		finv_table[ 608] = 36'b101000001010000010100000110010010111;
		finv_table[ 609] = 36'b101000001000011101110000110010010011;
		finv_table[ 610] = 36'b101000000110111001001100110010001111;
		finv_table[ 611] = 36'b101000000101010100101100110010001011;
		finv_table[ 612] = 36'b101000000011110000010110110010000111;
		finv_table[ 613] = 36'b101000000010001100001000110010000011;
		finv_table[ 614] = 36'b101000000000101000000000110001111111;
		finv_table[ 615] = 36'b100111111111000100000010110001111011;
		finv_table[ 616] = 36'b100111111101100000001010110001110111;
		finv_table[ 617] = 36'b100111111011111100011010110001110011;
		finv_table[ 618] = 36'b100111111010011000110010110001110000;
		finv_table[ 619] = 36'b100111111000110101010010110001101100;
		finv_table[ 620] = 36'b100111110111010001111010110001101000;
		finv_table[ 621] = 36'b100111110101101110101000110001100100;
		finv_table[ 622] = 36'b100111110100001011100000110001100000;
		finv_table[ 623] = 36'b100111110010101000011110110001011100;
		finv_table[ 624] = 36'b100111110001000101100100110001011000;
		finv_table[ 625] = 36'b100111101111100010110010110001010101;
		finv_table[ 626] = 36'b100111101110000000001010110001010001;
		finv_table[ 627] = 36'b100111101100011101100110110001001101;
		finv_table[ 628] = 36'b100111101010111011001100110001001001;
		finv_table[ 629] = 36'b100111101001011000111000110001000101;
		finv_table[ 630] = 36'b100111100111110110101110110001000010;
		finv_table[ 631] = 36'b100111100110010100101010110000111110;
		finv_table[ 632] = 36'b100111100100110010101100110000111010;
		finv_table[ 633] = 36'b100111100011010000111000110000110110;
		finv_table[ 634] = 36'b100111100001101111001010110000110010;
		finv_table[ 635] = 36'b100111100000001101100100110000101111;
		finv_table[ 636] = 36'b100111011110101100000110110000101011;
		finv_table[ 637] = 36'b100111011101001010110000110000100111;
		finv_table[ 638] = 36'b100111011011101001100000110000100011;
		finv_table[ 639] = 36'b100111011010001000011000110000100000;
		finv_table[ 640] = 36'b100111011000100111011000110000011100;
		finv_table[ 641] = 36'b100111010111000110011110110000011000;
		finv_table[ 642] = 36'b100111010101100101101100110000010100;
		finv_table[ 643] = 36'b100111010100000101000010110000010001;
		finv_table[ 644] = 36'b100111010010100100100010110000001101;
		finv_table[ 645] = 36'b100111010001000100000110110000001001;
		finv_table[ 646] = 36'b100111001111100011110010110000000110;
		finv_table[ 647] = 36'b100111001110000011100110110000000010;
		finv_table[ 648] = 36'b100111001100100011100000101111111110;
		finv_table[ 649] = 36'b100111001011000011100100101111111011;
		finv_table[ 650] = 36'b100111001001100011101110101111110111;
		finv_table[ 651] = 36'b100111001000000011111110101111110011;
		finv_table[ 652] = 36'b100111000110100100010110101111110000;
		finv_table[ 653] = 36'b100111000101000100110110101111101100;
		finv_table[ 654] = 36'b100111000011100101011100101111101000;
		finv_table[ 655] = 36'b100111000010000110001010101111100101;
		finv_table[ 656] = 36'b100111000000100111000000101111100001;
		finv_table[ 657] = 36'b100110111111000111111100101111011110;
		finv_table[ 658] = 36'b100110111101101001000000101111011010;
		finv_table[ 659] = 36'b100110111100001010001100101111010110;
		finv_table[ 660] = 36'b100110111010101011011110101111010011;
		finv_table[ 661] = 36'b100110111001001100111000101111001111;
		finv_table[ 662] = 36'b100110110111101110011000101111001100;
		finv_table[ 663] = 36'b100110110110010000000000101111001000;
		finv_table[ 664] = 36'b100110110100110001101110101111000100;
		finv_table[ 665] = 36'b100110110011010011100110101111000001;
		finv_table[ 666] = 36'b100110110001110101100010101110111101;
		finv_table[ 667] = 36'b100110110000010111100110101110111010;
		finv_table[ 668] = 36'b100110101110111001110010101110110110;
		finv_table[ 669] = 36'b100110101101011100000110101110110011;
		finv_table[ 670] = 36'b100110101011111110100000101110101111;
		finv_table[ 671] = 36'b100110101010100001000000101110101100;
		finv_table[ 672] = 36'b100110101001000011101000101110101000;
		finv_table[ 673] = 36'b100110100111100110010110101110100101;
		finv_table[ 674] = 36'b100110100110001001001100101110100001;
		finv_table[ 675] = 36'b100110100100101100001000101110011110;
		finv_table[ 676] = 36'b100110100011001111001100101110011010;
		finv_table[ 677] = 36'b100110100001110010010110101110010111;
		finv_table[ 678] = 36'b100110100000010101101010101110010011;
		finv_table[ 679] = 36'b100110011110111001000010101110010000;
		finv_table[ 680] = 36'b100110011101011100100010101110001100;
		finv_table[ 681] = 36'b100110011100000000001010101110001001;
		finv_table[ 682] = 36'b100110011010100011111000101110000101;
		finv_table[ 683] = 36'b100110011001000111101100101110000010;
		finv_table[ 684] = 36'b100110010111101011100110101101111110;
		finv_table[ 685] = 36'b100110010110001111101010101101111011;
		finv_table[ 686] = 36'b100110010100110011110010101101110111;
		finv_table[ 687] = 36'b100110010011011000000010101101110100;
		finv_table[ 688] = 36'b100110010001111100011000101101110001;
		finv_table[ 689] = 36'b100110010000100000111000101101101101;
		finv_table[ 690] = 36'b100110001111000101011100101101101010;
		finv_table[ 691] = 36'b100110001101101010001000101101100110;
		finv_table[ 692] = 36'b100110001100001110111010101101100011;
		finv_table[ 693] = 36'b100110001010110011110100101101100000;
		finv_table[ 694] = 36'b100110001001011000110100101101011100;
		finv_table[ 695] = 36'b100110000111111101111010101101011001;
		finv_table[ 696] = 36'b100110000110100011001000101101010101;
		finv_table[ 697] = 36'b100110000101001000011100101101010010;
		finv_table[ 698] = 36'b100110000011101101110110101101001111;
		finv_table[ 699] = 36'b100110000010010011011000101101001011;
		finv_table[ 700] = 36'b100110000000111001000000101101001000;
		finv_table[ 701] = 36'b100101111111011110110000101101000101;
		finv_table[ 702] = 36'b100101111110000100100110101101000001;
		finv_table[ 703] = 36'b100101111100101010100010101100111110;
		finv_table[ 704] = 36'b100101111011010000100100101100111011;
		finv_table[ 705] = 36'b100101111001110110110000101100110111;
		finv_table[ 706] = 36'b100101111000011101000000101100110100;
		finv_table[ 707] = 36'b100101110111000011010110101100110001;
		finv_table[ 708] = 36'b100101110101101001110100101100101101;
		finv_table[ 709] = 36'b100101110100010000011000101100101010;
		finv_table[ 710] = 36'b100101110010110111000010101100100111;
		finv_table[ 711] = 36'b100101110001011101110110101100100011;
		finv_table[ 712] = 36'b100101110000000100101110101100100000;
		finv_table[ 713] = 36'b100101101110101011101100101100011101;
		finv_table[ 714] = 36'b100101101101010010110010101100011010;
		finv_table[ 715] = 36'b100101101011111001111100101100010110;
		finv_table[ 716] = 36'b100101101010100001010000101100010011;
		finv_table[ 717] = 36'b100101101001001000101000101100010000;
		finv_table[ 718] = 36'b100101100111110000000110101100001101;
		finv_table[ 719] = 36'b100101100110010111101110101100001001;
		finv_table[ 720] = 36'b100101100100111111011010101100000110;
		finv_table[ 721] = 36'b100101100011100111001100101100000011;
		finv_table[ 722] = 36'b100101100010001111000110101100000000;
		finv_table[ 723] = 36'b100101100000110111000110101011111100;
		finv_table[ 724] = 36'b100101011111011111001100101011111001;
		finv_table[ 725] = 36'b100101011110000111011000101011110110;
		finv_table[ 726] = 36'b100101011100101111101010101011110011;
		finv_table[ 727] = 36'b100101011011011000000110101011110000;
		finv_table[ 728] = 36'b100101011010000000100100101011101100;
		finv_table[ 729] = 36'b100101011000101001001100101011101001;
		finv_table[ 730] = 36'b100101010111010001111000101011100110;
		finv_table[ 731] = 36'b100101010101111010101010101011100011;
		finv_table[ 732] = 36'b100101010100100011100100101011100000;
		finv_table[ 733] = 36'b100101010011001100100100101011011100;
		finv_table[ 734] = 36'b100101010001110101101010101011011001;
		finv_table[ 735] = 36'b100101010000011110110110101011010110;
		finv_table[ 736] = 36'b100101001111001000001010101011010011;
		finv_table[ 737] = 36'b100101001101110001100010101011010000;
		finv_table[ 738] = 36'b100101001100011011000010101011001101;
		finv_table[ 739] = 36'b100101001011000100100110101011001010;
		finv_table[ 740] = 36'b100101001001101110010010101011000110;
		finv_table[ 741] = 36'b100101001000011000000100101011000011;
		finv_table[ 742] = 36'b100101000111000001111100101011000000;
		finv_table[ 743] = 36'b100101000101101011111100101010111101;
		finv_table[ 744] = 36'b100101000100010110000000101010111010;
		finv_table[ 745] = 36'b100101000011000000001100101010110111;
		finv_table[ 746] = 36'b100101000001101010011100101010110100;
		finv_table[ 747] = 36'b100101000000010100110010101010110001;
		finv_table[ 748] = 36'b100100111110111111010010101010101110;
		finv_table[ 749] = 36'b100100111101101001110110101010101011;
		finv_table[ 750] = 36'b100100111100010100011110101010100111;
		finv_table[ 751] = 36'b100100111010111111001110101010100100;
		finv_table[ 752] = 36'b100100111001101010000110101010100001;
		finv_table[ 753] = 36'b100100111000010101000010101010011110;
		finv_table[ 754] = 36'b100100110111000000000100101010011011;
		finv_table[ 755] = 36'b100100110101101011001100101010011000;
		finv_table[ 756] = 36'b100100110100010110011100101010010101;
		finv_table[ 757] = 36'b100100110011000001110000101010010010;
		finv_table[ 758] = 36'b100100110001101101001100101010001111;
		finv_table[ 759] = 36'b100100110000011000101100101010001100;
		finv_table[ 760] = 36'b100100101111000100010100101010001001;
		finv_table[ 761] = 36'b100100101101110000000000101010000110;
		finv_table[ 762] = 36'b100100101100011011110100101010000011;
		finv_table[ 763] = 36'b100100101011000111101100101010000000;
		finv_table[ 764] = 36'b100100101001110011101100101001111101;
		finv_table[ 765] = 36'b100100101000011111110000101001111010;
		finv_table[ 766] = 36'b100100100111001011111100101001110111;
		finv_table[ 767] = 36'b100100100101111000001100101001110100;
		finv_table[ 768] = 36'b100100100100100100100100101001110001;
		finv_table[ 769] = 36'b100100100011010001000010101001101110;
		finv_table[ 770] = 36'b100100100001111101100100101001101011;
		finv_table[ 771] = 36'b100100100000101010001110101001101000;
		finv_table[ 772] = 36'b100100011111010110111100101001100101;
		finv_table[ 773] = 36'b100100011110000011110000101001100010;
		finv_table[ 774] = 36'b100100011100110000101100101001011111;
		finv_table[ 775] = 36'b100100011011011101101100101001011100;
		finv_table[ 776] = 36'b100100011010001010110100101001011001;
		finv_table[ 777] = 36'b100100011000111000000000101001010110;
		finv_table[ 778] = 36'b100100010111100101010010101001010011;
		finv_table[ 779] = 36'b100100010110010010101010101001010000;
		finv_table[ 780] = 36'b100100010101000000001000101001001110;
		finv_table[ 781] = 36'b100100010011101101101100101001001011;
		finv_table[ 782] = 36'b100100010010011011010110101001001000;
		finv_table[ 783] = 36'b100100010001001001001000101001000101;
		finv_table[ 784] = 36'b100100001111110110111100101001000010;
		finv_table[ 785] = 36'b100100001110100100111000101000111111;
		finv_table[ 786] = 36'b100100001101010010111000101000111100;
		finv_table[ 787] = 36'b100100001100000001000000101000111001;
		finv_table[ 788] = 36'b100100001010101111001100101000110110;
		finv_table[ 789] = 36'b100100001001011101011110101000110011;
		finv_table[ 790] = 36'b100100001000001011110110101000110001;
		finv_table[ 791] = 36'b100100000110111010010100101000101110;
		finv_table[ 792] = 36'b100100000101101000110110101000101011;
		finv_table[ 793] = 36'b100100000100010111100010101000101000;
		finv_table[ 794] = 36'b100100000011000110010010101000100101;
		finv_table[ 795] = 36'b100100000001110101000110101000100010;
		finv_table[ 796] = 36'b100100000000100100000000101000011111;
		finv_table[ 797] = 36'b100011111111010011000000101000011100;
		finv_table[ 798] = 36'b100011111110000010000110101000011010;
		finv_table[ 799] = 36'b100011111100110001010100101000010111;
		finv_table[ 800] = 36'b100011111011100000100100101000010100;
		finv_table[ 801] = 36'b100011111010001111111010101000010001;
		finv_table[ 802] = 36'b100011111000111111010110101000001110;
		finv_table[ 803] = 36'b100011110111101110111010101000001100;
		finv_table[ 804] = 36'b100011110110011110100010101000001001;
		finv_table[ 805] = 36'b100011110101001110001110101000000110;
		finv_table[ 806] = 36'b100011110011111110000010101000000011;
		finv_table[ 807] = 36'b100011110010101101111010101000000000;
		finv_table[ 808] = 36'b100011110001011101111010100111111110;
		finv_table[ 809] = 36'b100011110000001101111110100111111011;
		finv_table[ 810] = 36'b100011101110111110000110100111111000;
		finv_table[ 811] = 36'b100011101101101110010110100111110101;
		finv_table[ 812] = 36'b100011101100011110101010100111110010;
		finv_table[ 813] = 36'b100011101011001111000100100111110000;
		finv_table[ 814] = 36'b100011101001111111100100100111101101;
		finv_table[ 815] = 36'b100011101000110000001010100111101010;
		finv_table[ 816] = 36'b100011100111100000110110100111100111;
		finv_table[ 817] = 36'b100011100110010001100100100111100101;
		finv_table[ 818] = 36'b100011100101000010011100100111100010;
		finv_table[ 819] = 36'b100011100011110011011000100111011111;
		finv_table[ 820] = 36'b100011100010100100010110100111011100;
		finv_table[ 821] = 36'b100011100001010101011110100111011010;
		finv_table[ 822] = 36'b100011100000000110101010100111010111;
		finv_table[ 823] = 36'b100011011110110111111010100111010100;
		finv_table[ 824] = 36'b100011011101101001010010100111010001;
		finv_table[ 825] = 36'b100011011100011010101100100111001111;
		finv_table[ 826] = 36'b100011011011001100010000100111001100;
		finv_table[ 827] = 36'b100011011001111101110110100111001001;
		finv_table[ 828] = 36'b100011011000101111100010100111000111;
		finv_table[ 829] = 36'b100011010111100001010100100111000100;
		finv_table[ 830] = 36'b100011010110010011001100100111000001;
		finv_table[ 831] = 36'b100011010101000101001000100110111110;
		finv_table[ 832] = 36'b100011010011110111001010100110111100;
		finv_table[ 833] = 36'b100011010010101001010010100110111001;
		finv_table[ 834] = 36'b100011010001011011011110100110110110;
		finv_table[ 835] = 36'b100011010000001101110000100110110100;
		finv_table[ 836] = 36'b100011001111000000001000100110110001;
		finv_table[ 837] = 36'b100011001101110010100100100110101110;
		finv_table[ 838] = 36'b100011001100100101001000100110101100;
		finv_table[ 839] = 36'b100011001011010111110000100110101001;
		finv_table[ 840] = 36'b100011001010001010011010100110100110;
		finv_table[ 841] = 36'b100011001000111101001110100110100100;
		finv_table[ 842] = 36'b100011000111110000000110100110100001;
		finv_table[ 843] = 36'b100011000110100011000000100110011111;
		finv_table[ 844] = 36'b100011000101010110000100100110011100;
		finv_table[ 845] = 36'b100011000100001001001100100110011001;
		finv_table[ 846] = 36'b100011000010111100010110100110010111;
		finv_table[ 847] = 36'b100011000001101111101010100110010100;
		finv_table[ 848] = 36'b100011000000100011000000100110010001;
		finv_table[ 849] = 36'b100010111111010110011110100110001111;
		finv_table[ 850] = 36'b100010111110001001111110100110001100;
		finv_table[ 851] = 36'b100010111100111101100100100110001010;
		finv_table[ 852] = 36'b100010111011110001010010100110000111;
		finv_table[ 853] = 36'b100010111010100101000000100110000100;
		finv_table[ 854] = 36'b100010111001011000111000100110000010;
		finv_table[ 855] = 36'b100010111000001100110100100101111111;
		finv_table[ 856] = 36'b100010110111000000110100100101111101;
		finv_table[ 857] = 36'b100010110101110100111010100101111010;
		finv_table[ 858] = 36'b100010110100101001000100100101110111;
		finv_table[ 859] = 36'b100010110011011101010100100101110101;
		finv_table[ 860] = 36'b100010110010010001101010100101110010;
		finv_table[ 861] = 36'b100010110001000110000100100101110000;
		finv_table[ 862] = 36'b100010101111111010100100100101101101;
		finv_table[ 863] = 36'b100010101110101111001000100101101011;
		finv_table[ 864] = 36'b100010101101100011110010100101101000;
		finv_table[ 865] = 36'b100010101100011000100010100101100110;
		finv_table[ 866] = 36'b100010101011001101010110100101100011;
		finv_table[ 867] = 36'b100010101010000010001110100101100000;
		finv_table[ 868] = 36'b100010101000110111001100100101011110;
		finv_table[ 869] = 36'b100010100111101100010000100101011011;
		finv_table[ 870] = 36'b100010100110100001011010100101011001;
		finv_table[ 871] = 36'b100010100101010110100110100101010110;
		finv_table[ 872] = 36'b100010100100001011111000100101010100;
		finv_table[ 873] = 36'b100010100011000001010000100101010001;
		finv_table[ 874] = 36'b100010100001110110101100100101001111;
		finv_table[ 875] = 36'b100010100000101100001110100101001100;
		finv_table[ 876] = 36'b100010011111100001110100100101001010;
		finv_table[ 877] = 36'b100010011110010111100000100101000111;
		finv_table[ 878] = 36'b100010011101001101010000100101000101;
		finv_table[ 879] = 36'b100010011100000011000110100101000010;
		finv_table[ 880] = 36'b100010011010111001000000100101000000;
		finv_table[ 881] = 36'b100010011001101111000000100100111101;
		finv_table[ 882] = 36'b100010011000100101000100100100111011;
		finv_table[ 883] = 36'b100010010111011011001110100100111000;
		finv_table[ 884] = 36'b100010010110010001011100100100110110;
		finv_table[ 885] = 36'b100010010101000111110000100100110011;
		finv_table[ 886] = 36'b100010010011111110001000100100110001;
		finv_table[ 887] = 36'b100010010010110100100100100100101110;
		finv_table[ 888] = 36'b100010010001101011000110100100101100;
		finv_table[ 889] = 36'b100010010000100001101110100100101010;
		finv_table[ 890] = 36'b100010001111011000011010100100100111;
		finv_table[ 891] = 36'b100010001110001111001010100100100101;
		finv_table[ 892] = 36'b100010001101000110000000100100100010;
		finv_table[ 893] = 36'b100010001011111100111010100100100000;
		finv_table[ 894] = 36'b100010001010110011111010100100011101;
		finv_table[ 895] = 36'b100010001001101010111110100100011011;
		finv_table[ 896] = 36'b100010001000100010001000100100011000;
		finv_table[ 897] = 36'b100010000111011001010110100100010110;
		finv_table[ 898] = 36'b100010000110010000101010100100010100;
		finv_table[ 899] = 36'b100010000101001000000010100100010001;
		finv_table[ 900] = 36'b100010000011111111011110100100001111;
		finv_table[ 901] = 36'b100010000010110110111110100100001100;
		finv_table[ 902] = 36'b100010000001101110100110100100001010;
		finv_table[ 903] = 36'b100010000000100110010000100100001000;
		finv_table[ 904] = 36'b100001111111011110000000100100000101;
		finv_table[ 905] = 36'b100001111110010101110100100100000011;
		finv_table[ 906] = 36'b100001111101001101101110100100000000;
		finv_table[ 907] = 36'b100001111100000101101100100011111110;
		finv_table[ 908] = 36'b100001111010111101110000100011111100;
		finv_table[ 909] = 36'b100001111001110101111000100011111001;
		finv_table[ 910] = 36'b100001111000101110000100100011110111;
		finv_table[ 911] = 36'b100001110111100110010100100011110100;
		finv_table[ 912] = 36'b100001110110011110101010100011110010;
		finv_table[ 913] = 36'b100001110101010111000110100011110000;
		finv_table[ 914] = 36'b100001110100001111100110100011101101;
		finv_table[ 915] = 36'b100001110011001000001010100011101011;
		finv_table[ 916] = 36'b100001110010000000110100100011101001;
		finv_table[ 917] = 36'b100001110000111001100000100011100110;
		finv_table[ 918] = 36'b100001101111110010010010100011100100;
		finv_table[ 919] = 36'b100001101110101011001010100011100010;
		finv_table[ 920] = 36'b100001101101100100000110100011011111;
		finv_table[ 921] = 36'b100001101100011101000110100011011101;
		finv_table[ 922] = 36'b100001101011010110001100100011011011;
		finv_table[ 923] = 36'b100001101010001111010100100011011000;
		finv_table[ 924] = 36'b100001101001001000100010100011010110;
		finv_table[ 925] = 36'b100001101000000001110110100011010100;
		finv_table[ 926] = 36'b100001100110111011001110100011010001;
		finv_table[ 927] = 36'b100001100101110100101010100011001111;
		finv_table[ 928] = 36'b100001100100101110001010100011001101;
		finv_table[ 929] = 36'b100001100011100111101110100011001010;
		finv_table[ 930] = 36'b100001100010100001011010100011001000;
		finv_table[ 931] = 36'b100001100001011011001000100011000110;
		finv_table[ 932] = 36'b100001100000010100111100100011000100;
		finv_table[ 933] = 36'b100001011111001110110100100011000001;
		finv_table[ 934] = 36'b100001011110001000110010100010111111;
		finv_table[ 935] = 36'b100001011101000010110010100010111101;
		finv_table[ 936] = 36'b100001011011111100110110100010111010;
		finv_table[ 937] = 36'b100001011010110111000000100010111000;
		finv_table[ 938] = 36'b100001011001110001010000100010110110;
		finv_table[ 939] = 36'b100001011000101011100100100010110100;
		finv_table[ 940] = 36'b100001010111100101111100100010110001;
		finv_table[ 941] = 36'b100001010110100000011000100010101111;
		finv_table[ 942] = 36'b100001010101011010111010100010101101;
		finv_table[ 943] = 36'b100001010100010101011110100010101011;
		finv_table[ 944] = 36'b100001010011010000001000100010101000;
		finv_table[ 945] = 36'b100001010010001010110110100010100110;
		finv_table[ 946] = 36'b100001010001000101101010100010100100;
		finv_table[ 947] = 36'b100001010000000000100000100010100010;
		finv_table[ 948] = 36'b100001001110111011011110100010011111;
		finv_table[ 949] = 36'b100001001101110110011110100010011101;
		finv_table[ 950] = 36'b100001001100110001100100100010011011;
		finv_table[ 951] = 36'b100001001011101100101010100010011001;
		finv_table[ 952] = 36'b100001001010100111111000100010010110;
		finv_table[ 953] = 36'b100001001001100011001100100010010100;
		finv_table[ 954] = 36'b100001001000011110100010100010010010;
		finv_table[ 955] = 36'b100001000111011001111110100010010000;
		finv_table[ 956] = 36'b100001000110010101011110100010001101;
		finv_table[ 957] = 36'b100001000101010001000010100010001011;
		finv_table[ 958] = 36'b100001000100001100101010100010001001;
		finv_table[ 959] = 36'b100001000011001000011000100010000111;
		finv_table[ 960] = 36'b100001000010000100001000100010000101;
		finv_table[ 961] = 36'b100001000000111111111100100010000010;
		finv_table[ 962] = 36'b100000111111111011111000100010000000;
		finv_table[ 963] = 36'b100000111110110111110110100001111110;
		finv_table[ 964] = 36'b100000111101110011111000100001111100;
		finv_table[ 965] = 36'b100000111100110000000000100001111010;
		finv_table[ 966] = 36'b100000111011101100001100100001111000;
		finv_table[ 967] = 36'b100000111010101000011100100001110101;
		finv_table[ 968] = 36'b100000111001100100110000100001110011;
		finv_table[ 969] = 36'b100000111000100001001010100001110001;
		finv_table[ 970] = 36'b100000110111011101100110100001101111;
		finv_table[ 971] = 36'b100000110110011010000110100001101101;
		finv_table[ 972] = 36'b100000110101010110101100100001101011;
		finv_table[ 973] = 36'b100000110100010011010110100001101000;
		finv_table[ 974] = 36'b100000110011010000000100100001100110;
		finv_table[ 975] = 36'b100000110010001100111000100001100100;
		finv_table[ 976] = 36'b100000110001001001101110100001100010;
		finv_table[ 977] = 36'b100000110000000110101010100001100000;
		finv_table[ 978] = 36'b100000101111000011101000100001011110;
		finv_table[ 979] = 36'b100000101110000000101100100001011011;
		finv_table[ 980] = 36'b100000101100111101110100100001011001;
		finv_table[ 981] = 36'b100000101011111011000010100001010111;
		finv_table[ 982] = 36'b100000101010111000010010100001010101;
		finv_table[ 983] = 36'b100000101001110101101000100001010011;
		finv_table[ 984] = 36'b100000101000110011000000100001010001;
		finv_table[ 985] = 36'b100000100111110000011100100001001111;
		finv_table[ 986] = 36'b100000100110101110000000100001001101;
		finv_table[ 987] = 36'b100000100101101011100100100001001010;
		finv_table[ 988] = 36'b100000100100101001001110100001001000;
		finv_table[ 989] = 36'b100000100011100110111100100001000110;
		finv_table[ 990] = 36'b100000100010100100101110100001000100;
		finv_table[ 991] = 36'b100000100001100010100110100001000010;
		finv_table[ 992] = 36'b100000100000100000100000100001000000;
		finv_table[ 993] = 36'b100000011111011110100000100000111110;
		finv_table[ 994] = 36'b100000011110011100100010100000111100;
		finv_table[ 995] = 36'b100000011101011010101010100000111010;
		finv_table[ 996] = 36'b100000011100011000110110100000111000;
		finv_table[ 997] = 36'b100000011011010111000100100000110110;
		finv_table[ 998] = 36'b100000011010010101011000100000110011;
		finv_table[ 999] = 36'b100000011001010011110010100000110001;
		finv_table[1000] = 36'b100000011000010010001110100000101111;
		finv_table[1001] = 36'b100000010111010000101110100000101101;
		finv_table[1002] = 36'b100000010110001111010010100000101011;
		finv_table[1003] = 36'b100000010101001101111100100000101001;
		finv_table[1004] = 36'b100000010100001100101000100000100111;
		finv_table[1005] = 36'b100000010011001011011010100000100101;
		finv_table[1006] = 36'b100000010010001010001110100000100011;
		finv_table[1007] = 36'b100000010001001001001000100000100001;
		finv_table[1008] = 36'b100000010000001000000100100000011111;
		finv_table[1009] = 36'b100000001111000111000100100000011101;
		finv_table[1010] = 36'b100000001110000110001100100000011011;
		finv_table[1011] = 36'b100000001101000101010010100000011001;
		finv_table[1012] = 36'b100000001100000100100010100000010111;
		finv_table[1013] = 36'b100000001011000011110010100000010101;
		finv_table[1014] = 36'b100000001010000011001000100000010011;
		finv_table[1015] = 36'b100000001001000010100010100000010001;
		finv_table[1016] = 36'b100000001000000010000010100000001111;
		finv_table[1017] = 36'b100000000111000001100010100000001101;
		finv_table[1018] = 36'b100000000110000001001000100000001011;
		finv_table[1019] = 36'b100000000101000000110010100000001001;
		finv_table[1020] = 36'b100000000100000000100000100000000111;
		finv_table[1021] = 36'b100000000011000000010010100000000101;
		finv_table[1022] = 36'b100000000010000000001000100000000011;
		finv_table[1023] = 36'b100000000001000000000010100000000001;
	end
endmodule

`default_nettype wire