`default_nettype none
module sqrt (
	input wire [31:0]  x,
  output wire [31:0] y,
  //output wire        ovf,
  input wire       clk,
  input wire       rstn
);
	wire     	 	sign = x[31];
	wire [ 7:0] exp_x = x[30:23];
	wire [22:0] frac_x = x[22:0];
	wire [ 7:0] exp_x_unbiased = exp_x - 8'd127;

	wire [ 9:0] addr = {exp_x_unbiased[0],x[22:14]};
	wire [13:0] dx = x[13:0];
	wire [35:0] dout;
	sqrt_table sqrt_table1(addr, dout, clk, rstn);

	wire [22:0] constant = dout[35:13];
	wire [12:0] gradient = dout[12:0];
	wire [26:0] dy_calc = gradient * dx;
	wire [22:0] frac_y = constant + dy_calc[26:4];

	wire [ 7:0] exp_y_unbiased = exp_x_unbiased >> 1;
	wire [ 7:0] exp_y = exp_y_unbiased + 8'd127;

	assign y = {sign , exp_y, frac_y};
endmodule

module sqrt_table (
	input		wire [ 9:0]	addr,
	output	reg  [35:0] dout,
	input 	wire 				clk,
	input 	wire 				rstn
);
	(*ram_style = "BLOCK"*) logic [35:0] sqrt_table [1023:0];
	always @(posedge clk) begin
		dout <= sqrt_table[addr];
	end
	initial begin
		sqrt_table[   0] = 36'b000000000000000000000000111111111110;
		sqrt_table[   1] = 36'b000000000011111111111000111111111010;
		sqrt_table[   2] = 36'b000000000111111111100000111111110110;
		sqrt_table[   3] = 36'b000000001011111110111000111111110010;
		sqrt_table[   4] = 36'b000000001111111110000000111111101110;
		sqrt_table[   5] = 36'b000000010011111100111000111111101010;
		sqrt_table[   6] = 36'b000000010111111011100100111111100110;
		sqrt_table[   7] = 36'b000000011011111001111100111111100010;
		sqrt_table[   8] = 36'b000000011111111000000100111111011110;
		sqrt_table[   9] = 36'b000000100011110110000000111111011010;
		sqrt_table[  10] = 36'b000000100111110011101000111111010110;
		sqrt_table[  11] = 36'b000000101011110001000010111111010011;
		sqrt_table[  12] = 36'b000000101111101110010000111111001110;
		sqrt_table[  13] = 36'b000000110011101011001000111111001011;
		sqrt_table[  14] = 36'b000000110111100111110110111111000111;
		sqrt_table[  15] = 36'b000000111011100100010000111111000011;
		sqrt_table[  16] = 36'b000000111111100000100000111110111111;
		sqrt_table[  17] = 36'b000001000011011100011100111110111011;
		sqrt_table[  18] = 36'b000001000111011000001100111110111000;
		sqrt_table[  19] = 36'b000001001011010011101100111110110100;
		sqrt_table[  20] = 36'b000001001111001111000000111110110000;
		sqrt_table[  21] = 36'b000001010011001001111110111110101101;
		sqrt_table[  22] = 36'b000001010111000100110100111110101000;
		sqrt_table[  23] = 36'b000001011010111111010110111110100101;
		sqrt_table[  24] = 36'b000001011110111001101000111110100001;
		sqrt_table[  25] = 36'b000001100010110011110000111110011110;
		sqrt_table[  26] = 36'b000001100110101101100100111110011001;
		sqrt_table[  27] = 36'b000001101010100111001100111110010110;
		sqrt_table[  28] = 36'b000001101110100000101000111110010010;
		sqrt_table[  29] = 36'b000001110010011001110010111110001111;
		sqrt_table[  30] = 36'b000001110110010010101110111110001011;
		sqrt_table[  31] = 36'b000001111010001011011000111110000111;
		sqrt_table[  32] = 36'b000001111110000011111000111110000100;
		sqrt_table[  33] = 36'b000010000001111100001000111110000000;
		sqrt_table[  34] = 36'b000010000101110100000110111101111101;
		sqrt_table[  35] = 36'b000010001001101011111010111101111001;
		sqrt_table[  36] = 36'b000010001101100011011110111101110101;
		sqrt_table[  37] = 36'b000010010001011010110100111101110010;
		sqrt_table[  38] = 36'b000010010101010001111100111101101110;
		sqrt_table[  39] = 36'b000010011001001000110100111101101010;
		sqrt_table[  40] = 36'b000010011100111111011110111101100111;
		sqrt_table[  41] = 36'b000010100000110101111000111101100011;
		sqrt_table[  42] = 36'b000010100100101100001000111101100000;
		sqrt_table[  43] = 36'b000010101000100010001000111101011100;
		sqrt_table[  44] = 36'b000010101100010111111010111101011001;
		sqrt_table[  45] = 36'b000010110000001101011110111101010101;
		sqrt_table[  46] = 36'b000010110100000010110000111101010010;
		sqrt_table[  47] = 36'b000010110111110111111000111101001110;
		sqrt_table[  48] = 36'b000010111011101100110010111101001011;
		sqrt_table[  49] = 36'b000010111111100001011110111101000111;
		sqrt_table[  50] = 36'b000011000011010101111000111101000100;
		sqrt_table[  51] = 36'b000011000111001010001000111101000000;
		sqrt_table[  52] = 36'b000011001010111110001100111100111100;
		sqrt_table[  53] = 36'b000011001110110001111100111100111001;
		sqrt_table[  54] = 36'b000011010010100101100100111100110110;
		sqrt_table[  55] = 36'b000011010110011000111100111100110010;
		sqrt_table[  56] = 36'b000011011010001100000100111100101111;
		sqrt_table[  57] = 36'b000011011101111111000000111100101011;
		sqrt_table[  58] = 36'b000011100001110001110000111100101000;
		sqrt_table[  59] = 36'b000011100101100100010010111100100101;
		sqrt_table[  60] = 36'b000011101001010110100100111100100001;
		sqrt_table[  61] = 36'b000011101101001000101100111100011110;
		sqrt_table[  62] = 36'b000011110000111010100110111100011011;
		sqrt_table[  63] = 36'b000011110100101100010010111100010111;
		sqrt_table[  64] = 36'b000011111000011101101100111100010100;
		sqrt_table[  65] = 36'b000011111100001111000000111100010000;
		sqrt_table[  66] = 36'b000100000000000000000000111100001101;
		sqrt_table[  67] = 36'b000100000011110000111000111100001010;
		sqrt_table[  68] = 36'b000100000111100001100000111100000110;
		sqrt_table[  69] = 36'b000100001011010001111000111100000011;
		sqrt_table[  70] = 36'b000100001111000010001000111100000000;
		sqrt_table[  71] = 36'b000100010010110010001000111011111100;
		sqrt_table[  72] = 36'b000100010110100001111100111011111001;
		sqrt_table[  73] = 36'b000100011010010001100000111011110110;
		sqrt_table[  74] = 36'b000100011110000000111010111011110011;
		sqrt_table[  75] = 36'b000100100001110000001000111011110000;
		sqrt_table[  76] = 36'b000100100101011111001000111011101100;
		sqrt_table[  77] = 36'b000100101001001101111010111011101001;
		sqrt_table[  78] = 36'b000100101100111100011100111011100110;
		sqrt_table[  79] = 36'b000100110000101010110110111011100011;
		sqrt_table[  80] = 36'b000100110100011001000000111011011111;
		sqrt_table[  81] = 36'b000100111000000111000000111011011100;
		sqrt_table[  82] = 36'b000100111011110100110010111011011001;
		sqrt_table[  83] = 36'b000100111111100010010100111011010110;
		sqrt_table[  84] = 36'b000101000011001111101110111011010011;
		sqrt_table[  85] = 36'b000101000110111100111000111011001111;
		sqrt_table[  86] = 36'b000101001010101001111000111011001100;
		sqrt_table[  87] = 36'b000101001110010110101000111011001001;
		sqrt_table[  88] = 36'b000101010010000011001110111011000110;
		sqrt_table[  89] = 36'b000101010101101111100110111011000011;
		sqrt_table[  90] = 36'b000101011001011011110010111011000000;
		sqrt_table[  91] = 36'b000101011101000111110100111010111100;
		sqrt_table[  92] = 36'b000101100000110011100100111010111001;
		sqrt_table[  93] = 36'b000101100100011111001100111010110110;
		sqrt_table[  94] = 36'b000101101000001010100100111010110011;
		sqrt_table[  95] = 36'b000101101011110101110100111010110000;
		sqrt_table[  96] = 36'b000101101111100000110110111010101101;
		sqrt_table[  97] = 36'b000101110011001011101000111010101010;
		sqrt_table[  98] = 36'b000101110110110110010010111010100111;
		sqrt_table[  99] = 36'b000101111010100000101100111010100100;
		sqrt_table[ 100] = 36'b000101111110001010111110111010100001;
		sqrt_table[ 101] = 36'b000110000001110101000000111010011110;
		sqrt_table[ 102] = 36'b000110000101011110111000111010011011;
		sqrt_table[ 103] = 36'b000110001001001000100100111010010111;
		sqrt_table[ 104] = 36'b000110001100110010000010111010010101;
		sqrt_table[ 105] = 36'b000110010000011011010100111010010001;
		sqrt_table[ 106] = 36'b000110010100000100011100111010001110;
		sqrt_table[ 107] = 36'b000110010111101101011000111010001100;
		sqrt_table[ 108] = 36'b000110011011010110001000111010001000;
		sqrt_table[ 109] = 36'b000110011110111110101000111010000110;
		sqrt_table[ 110] = 36'b000110100010100111000000111010000010;
		sqrt_table[ 111] = 36'b000110100110001111001000111001111111;
		sqrt_table[ 112] = 36'b000110101001110111001010111001111101;
		sqrt_table[ 113] = 36'b000110101101011110111100111001111010;
		sqrt_table[ 114] = 36'b000110110001000110100100111001110110;
		sqrt_table[ 115] = 36'b000110110100101110000000111001110100;
		sqrt_table[ 116] = 36'b000110111000010101001110111001110001;
		sqrt_table[ 117] = 36'b000110111011111100010100111001101110;
		sqrt_table[ 118] = 36'b000110111111100011001010111001101011;
		sqrt_table[ 119] = 36'b000111000011001001111000111001101000;
		sqrt_table[ 120] = 36'b000111000110110000010100111001100101;
		sqrt_table[ 121] = 36'b000111001010010110101100111001100010;
		sqrt_table[ 122] = 36'b000111001101111100110100111001011111;
		sqrt_table[ 123] = 36'b000111010001100010110100111001011100;
		sqrt_table[ 124] = 36'b000111010101001000100100111001011010;
		sqrt_table[ 125] = 36'b000111011000101110001100111001010110;
		sqrt_table[ 126] = 36'b000111011100010011101000111001010100;
		sqrt_table[ 127] = 36'b000111011111111000110110111001010001;
		sqrt_table[ 128] = 36'b000111100011011101111100111001001110;
		sqrt_table[ 129] = 36'b000111100111000010110000111001001011;
		sqrt_table[ 130] = 36'b000111101010100111100000111001001000;
		sqrt_table[ 131] = 36'b000111101110001100000000111001000101;
		sqrt_table[ 132] = 36'b000111110001110000011000111001000010;
		sqrt_table[ 133] = 36'b000111110101010100100100111001000000;
		sqrt_table[ 134] = 36'b000111111000111000100010111000111101;
		sqrt_table[ 135] = 36'b000111111100011100011000111000111010;
		sqrt_table[ 136] = 36'b001000000000000000000000111000110111;
		sqrt_table[ 137] = 36'b001000000011100011100000111000110100;
		sqrt_table[ 138] = 36'b001000000111000110110000111000110010;
		sqrt_table[ 139] = 36'b001000001010101001111010111000101111;
		sqrt_table[ 140] = 36'b001000001110001100110100111000101100;
		sqrt_table[ 141] = 36'b001000010001101111100100111000101001;
		sqrt_table[ 142] = 36'b001000010101010010001100111000100111;
		sqrt_table[ 143] = 36'b001000011000110100101000111000100100;
		sqrt_table[ 144] = 36'b001000011100010110111000111000100001;
		sqrt_table[ 145] = 36'b001000011111111000111100111000011110;
		sqrt_table[ 146] = 36'b001000100011011010110100111000011011;
		sqrt_table[ 147] = 36'b001000100110111100100110111000011001;
		sqrt_table[ 148] = 36'b001000101010011110001000111000010110;
		sqrt_table[ 149] = 36'b001000101101111111100000111000010011;
		sqrt_table[ 150] = 36'b001000110001100000110010111000010001;
		sqrt_table[ 151] = 36'b001000110101000001110100111000001110;
		sqrt_table[ 152] = 36'b001000111000100010101100111000001011;
		sqrt_table[ 153] = 36'b001000111100000011011100111000001000;
		sqrt_table[ 154] = 36'b001000111111100011111100111000000110;
		sqrt_table[ 155] = 36'b001001000011000100010100111000000011;
		sqrt_table[ 156] = 36'b001001000110100100100100111000000000;
		sqrt_table[ 157] = 36'b001001001010000100100100110111111110;
		sqrt_table[ 158] = 36'b001001001101100100011100110111111011;
		sqrt_table[ 159] = 36'b001001010001000100001100110111111000;
		sqrt_table[ 160] = 36'b001001010100100011101100110111110110;
		sqrt_table[ 161] = 36'b001001011000000011000110110111110011;
		sqrt_table[ 162] = 36'b001001011011100010010010110111110001;
		sqrt_table[ 163] = 36'b001001011111000001010100110111101110;
		sqrt_table[ 164] = 36'b001001100010100000001110110111101011;
		sqrt_table[ 165] = 36'b001001100101111110111010110111101001;
		sqrt_table[ 166] = 36'b001001101001011101011100110111100110;
		sqrt_table[ 167] = 36'b001001101100111011110100110111100011;
		sqrt_table[ 168] = 36'b001001110000011010000010110111100001;
		sqrt_table[ 169] = 36'b001001110011111000001000110111011110;
		sqrt_table[ 170] = 36'b001001110111010110000000110111011100;
		sqrt_table[ 171] = 36'b001001111010110011101110110111011001;
		sqrt_table[ 172] = 36'b001001111110010001010100110111010110;
		sqrt_table[ 173] = 36'b001010000001101110101100110111010100;
		sqrt_table[ 174] = 36'b001010000101001011111110110111010001;
		sqrt_table[ 175] = 36'b001010001000101001000010110111001111;
		sqrt_table[ 176] = 36'b001010001100000101111100110111001100;
		sqrt_table[ 177] = 36'b001010001111100010101100110111001001;
		sqrt_table[ 178] = 36'b001010010010111111010000110111000111;
		sqrt_table[ 179] = 36'b001010010110011011110000110111000100;
		sqrt_table[ 180] = 36'b001010011001111000000000110111000001;
		sqrt_table[ 181] = 36'b001010011101010100001000110110111111;
		sqrt_table[ 182] = 36'b001010100000110000000110110110111101;
		sqrt_table[ 183] = 36'b001010100100001011111100110110111010;
		sqrt_table[ 184] = 36'b001010100111100111100100110110110111;
		sqrt_table[ 185] = 36'b001010101011000011000000110110110101;
		sqrt_table[ 186] = 36'b001010101110011110011010110110110011;
		sqrt_table[ 187] = 36'b001010110001111001100100110110110000;
		sqrt_table[ 188] = 36'b001010110101010100100100110110101110;
		sqrt_table[ 189] = 36'b001010111000101111011100110110101011;
		sqrt_table[ 190] = 36'b001010111100001010001100110110101000;
		sqrt_table[ 191] = 36'b001010111111100100101100110110100110;
		sqrt_table[ 192] = 36'b001011000010111111000100110110100011;
		sqrt_table[ 193] = 36'b001011000110011001010100110110100001;
		sqrt_table[ 194] = 36'b001011001001110011011010110110011111;
		sqrt_table[ 195] = 36'b001011001101001101011000110110011100;
		sqrt_table[ 196] = 36'b001011010000100111001000110110011010;
		sqrt_table[ 197] = 36'b001011010100000000110000110110010111;
		sqrt_table[ 198] = 36'b001011010111011010001110110110010101;
		sqrt_table[ 199] = 36'b001011011010110011100100110110010010;
		sqrt_table[ 200] = 36'b001011011110001100101100110110010000;
		sqrt_table[ 201] = 36'b001011100001100101101100110110001101;
		sqrt_table[ 202] = 36'b001011100100111110100100110110001011;
		sqrt_table[ 203] = 36'b001011101000010111010100110110001000;
		sqrt_table[ 204] = 36'b001011101011101111110100110110000110;
		sqrt_table[ 205] = 36'b001011101111001000010000110110000100;
		sqrt_table[ 206] = 36'b001011110010100000100000110110000001;
		sqrt_table[ 207] = 36'b001011110101111000100110110101111111;
		sqrt_table[ 208] = 36'b001011111001010000100010110101111101;
		sqrt_table[ 209] = 36'b001011111100101000011000110101111010;
		sqrt_table[ 210] = 36'b001100000000000000000000110101111000;
		sqrt_table[ 211] = 36'b001100000011010111100000110101110110;
		sqrt_table[ 212] = 36'b001100000110101110111000110101110011;
		sqrt_table[ 213] = 36'b001100001010000110000110110101110001;
		sqrt_table[ 214] = 36'b001100001101011101001000110101101110;
		sqrt_table[ 215] = 36'b001100010000110100000100110101101100;
		sqrt_table[ 216] = 36'b001100010100001010110100110101101001;
		sqrt_table[ 217] = 36'b001100010111100001011000110101100111;
		sqrt_table[ 218] = 36'b001100011010110111111010110101100101;
		sqrt_table[ 219] = 36'b001100011110001110001110110101100011;
		sqrt_table[ 220] = 36'b001100100001100100011000110101100000;
		sqrt_table[ 221] = 36'b001100100100111010011100110101011110;
		sqrt_table[ 222] = 36'b001100101000010000010100110101011100;
		sqrt_table[ 223] = 36'b001100101011100110000000110101011001;
		sqrt_table[ 224] = 36'b001100101110111011101000110101010111;
		sqrt_table[ 225] = 36'b001100110010010001000100110101010101;
		sqrt_table[ 226] = 36'b001100110101100110011000110101010010;
		sqrt_table[ 227] = 36'b001100111000111011100010110101010000;
		sqrt_table[ 228] = 36'b001100111100010000100100110101001110;
		sqrt_table[ 229] = 36'b001100111111100101011000110101001011;
		sqrt_table[ 230] = 36'b001101000010111010001000110101001001;
		sqrt_table[ 231] = 36'b001101000110001110101110110101000111;
		sqrt_table[ 232] = 36'b001101001001100011001100110101000100;
		sqrt_table[ 233] = 36'b001101001100110111011100110101000010;
		sqrt_table[ 234] = 36'b001101010000001011101000110101000000;
		sqrt_table[ 235] = 36'b001101010011011111101000110100111101;
		sqrt_table[ 236] = 36'b001101010110110011100000110100111100;
		sqrt_table[ 237] = 36'b001101011010000111001110110100111001;
		sqrt_table[ 238] = 36'b001101011101011010110000110100110111;
		sqrt_table[ 239] = 36'b001101100000101110010000110100110101;
		sqrt_table[ 240] = 36'b001101100100000001100100110100110010;
		sqrt_table[ 241] = 36'b001101100111010100110000110100110000;
		sqrt_table[ 242] = 36'b001101101010100111110000110100101110;
		sqrt_table[ 243] = 36'b001101101101111010101000110100101100;
		sqrt_table[ 244] = 36'b001101110001001101011000110100101001;
		sqrt_table[ 245] = 36'b001101110100011111111100110100100111;
		sqrt_table[ 246] = 36'b001101110111110010011100110100100101;
		sqrt_table[ 247] = 36'b001101111011000100110010110100100011;
		sqrt_table[ 248] = 36'b001101111110010111000000110100100000;
		sqrt_table[ 249] = 36'b001110000001101001000000110100011110;
		sqrt_table[ 250] = 36'b001110000100111010111100110100011100;
		sqrt_table[ 251] = 36'b001110001000001100101100110100011010;
		sqrt_table[ 252] = 36'b001110001011011110010110110100011000;
		sqrt_table[ 253] = 36'b001110001110101111110100110100010101;
		sqrt_table[ 254] = 36'b001110010010000001001100110100010100;
		sqrt_table[ 255] = 36'b001110010101010010011100110100010001;
		sqrt_table[ 256] = 36'b001110011000100011100010110100001111;
		sqrt_table[ 257] = 36'b001110011011110100011110110100001101;
		sqrt_table[ 258] = 36'b001110011111000101010010110100001011;
		sqrt_table[ 259] = 36'b001110100010010101111110110100001001;
		sqrt_table[ 260] = 36'b001110100101100110100100110100000110;
		sqrt_table[ 261] = 36'b001110101000110110111100110100000100;
		sqrt_table[ 262] = 36'b001110101100000111010000110100000010;
		sqrt_table[ 263] = 36'b001110101111010111011000110100000000;
		sqrt_table[ 264] = 36'b001110110010100111011000110011111110;
		sqrt_table[ 265] = 36'b001110110101110111010000110011111100;
		sqrt_table[ 266] = 36'b001110111001000111000000110011111001;
		sqrt_table[ 267] = 36'b001110111100010110100100110011110111;
		sqrt_table[ 268] = 36'b001110111111100110000100110011110101;
		sqrt_table[ 269] = 36'b001111000010110101011000110011110011;
		sqrt_table[ 270] = 36'b001111000110000100101000110011110001;
		sqrt_table[ 271] = 36'b001111001001010011101110110011101111;
		sqrt_table[ 272] = 36'b001111001100100010101010110011101101;
		sqrt_table[ 273] = 36'b001111001111110001011110110011101011;
		sqrt_table[ 274] = 36'b001111010011000000001100110011101000;
		sqrt_table[ 275] = 36'b001111010110001110101100110011100111;
		sqrt_table[ 276] = 36'b001111011001011101001000110011100100;
		sqrt_table[ 277] = 36'b001111011100101011011100110011100010;
		sqrt_table[ 278] = 36'b001111011111111001100100110011100000;
		sqrt_table[ 279] = 36'b001111100011000111101000110011011110;
		sqrt_table[ 280] = 36'b001111100110010101100000110011011100;
		sqrt_table[ 281] = 36'b001111101001100011010000110011011010;
		sqrt_table[ 282] = 36'b001111101100110000111000110011011000;
		sqrt_table[ 283] = 36'b001111101111111110011010110011010110;
		sqrt_table[ 284] = 36'b001111110011001011110010110011010100;
		sqrt_table[ 285] = 36'b001111110110011001000010110011010010;
		sqrt_table[ 286] = 36'b001111111001100110001000110011001111;
		sqrt_table[ 287] = 36'b001111111100110011001000110011001110;
		sqrt_table[ 288] = 36'b010000000000000000000000110011001100;
		sqrt_table[ 289] = 36'b010000000011001100110000110011001001;
		sqrt_table[ 290] = 36'b010000000110011001010100110011000111;
		sqrt_table[ 291] = 36'b010000001001100101110100110011000110;
		sqrt_table[ 292] = 36'b010000001100110010001100110011000011;
		sqrt_table[ 293] = 36'b010000001111111110011000110011000001;
		sqrt_table[ 294] = 36'b010000010011001010100000110010111111;
		sqrt_table[ 295] = 36'b010000010110010110011100110010111101;
		sqrt_table[ 296] = 36'b010000011001100010010100110010111011;
		sqrt_table[ 297] = 36'b010000011100101110000000110010111001;
		sqrt_table[ 298] = 36'b010000011111111001101000110010110111;
		sqrt_table[ 299] = 36'b010000100011000101000100110010110101;
		sqrt_table[ 300] = 36'b010000100110010000011100110010110011;
		sqrt_table[ 301] = 36'b010000101001011011101000110010110001;
		sqrt_table[ 302] = 36'b010000101100100110110000110010101111;
		sqrt_table[ 303] = 36'b010000101111110001101100110010101101;
		sqrt_table[ 304] = 36'b010000110010111100100100110010101100;
		sqrt_table[ 305] = 36'b010000110110000111010100110010101001;
		sqrt_table[ 306] = 36'b010000111001010001111000110010100111;
		sqrt_table[ 307] = 36'b010000111100011100011000110010100101;
		sqrt_table[ 308] = 36'b010000111111100110101100110010100011;
		sqrt_table[ 309] = 36'b010001000010110000111100110010100001;
		sqrt_table[ 310] = 36'b010001000101111011000100110010100000;
		sqrt_table[ 311] = 36'b010001001001000101000000110010011101;
		sqrt_table[ 312] = 36'b010001001100001110111000110010011100;
		sqrt_table[ 313] = 36'b010001001111011000101000110010011001;
		sqrt_table[ 314] = 36'b010001010010100010010000110010011000;
		sqrt_table[ 315] = 36'b010001010101101011101110110010010110;
		sqrt_table[ 316] = 36'b010001011000110101000110110010010100;
		sqrt_table[ 317] = 36'b010001011011111110010110110010010010;
		sqrt_table[ 318] = 36'b010001011111000111011110110010010000;
		sqrt_table[ 319] = 36'b010001100010010000011110110010001110;
		sqrt_table[ 320] = 36'b010001100101011001011000110010001100;
		sqrt_table[ 321] = 36'b010001101000100010001000110010001010;
		sqrt_table[ 322] = 36'b010001101011101010110000110010001000;
		sqrt_table[ 323] = 36'b010001101110110011010100110010000110;
		sqrt_table[ 324] = 36'b010001110001111011101010110010000101;
		sqrt_table[ 325] = 36'b010001110101000100000000110010000010;
		sqrt_table[ 326] = 36'b010001111000001100001000110010000000;
		sqrt_table[ 327] = 36'b010001111011010100001010110001111111;
		sqrt_table[ 328] = 36'b010001111110011100001000110001111100;
		sqrt_table[ 329] = 36'b010010000001100011111010110001111011;
		sqrt_table[ 330] = 36'b010010000100101011100100110001111001;
		sqrt_table[ 331] = 36'b010010000111110011001010110001110111;
		sqrt_table[ 332] = 36'b010010001010111010100110110001110101;
		sqrt_table[ 333] = 36'b010010001110000001111000110001110011;
		sqrt_table[ 334] = 36'b010010010001001001001000110001110001;
		sqrt_table[ 335] = 36'b010010010100010000001110110001110000;
		sqrt_table[ 336] = 36'b010010010111010111001100110001101101;
		sqrt_table[ 337] = 36'b010010011010011110000100110001101100;
		sqrt_table[ 338] = 36'b010010011101100100110100110001101010;
		sqrt_table[ 339] = 36'b010010100000101011011100110001101000;
		sqrt_table[ 340] = 36'b010010100011110001111100110001100110;
		sqrt_table[ 341] = 36'b010010100110111000011000110001100100;
		sqrt_table[ 342] = 36'b010010101001111110101000110001100010;
		sqrt_table[ 343] = 36'b010010101101000100110100110001100000;
		sqrt_table[ 344] = 36'b010010110000001010110110110001011111;
		sqrt_table[ 345] = 36'b010010110011010000110010110001011101;
		sqrt_table[ 346] = 36'b010010110110010110100100110001011011;
		sqrt_table[ 347] = 36'b010010111001011100010010110001011001;
		sqrt_table[ 348] = 36'b010010111100100001110100110001010111;
		sqrt_table[ 349] = 36'b010010111111100111010100110001010110;
		sqrt_table[ 350] = 36'b010011000010101100101100110001010011;
		sqrt_table[ 351] = 36'b010011000101110001111100110001010010;
		sqrt_table[ 352] = 36'b010011001000110111000100110001010000;
		sqrt_table[ 353] = 36'b010011001011111100000100110001001110;
		sqrt_table[ 354] = 36'b010011001111000001000000110001001100;
		sqrt_table[ 355] = 36'b010011010010000101110000110001001010;
		sqrt_table[ 356] = 36'b010011010101001010011010110001001001;
		sqrt_table[ 357] = 36'b010011011000001110111110110001000111;
		sqrt_table[ 358] = 36'b010011011011010011011000110001000101;
		sqrt_table[ 359] = 36'b010011011110010111110000110001000011;
		sqrt_table[ 360] = 36'b010011100001011011111100110001000001;
		sqrt_table[ 361] = 36'b010011100100100000000100110001000000;
		sqrt_table[ 362] = 36'b010011100111100100000100110000111110;
		sqrt_table[ 363] = 36'b010011101010100111111100110000111100;
		sqrt_table[ 364] = 36'b010011101101101011110000110000111010;
		sqrt_table[ 365] = 36'b010011110000101111011000110000111001;
		sqrt_table[ 366] = 36'b010011110011110010111100110000110110;
		sqrt_table[ 367] = 36'b010011110110110110010100110000110101;
		sqrt_table[ 368] = 36'b010011111001111001101100110000110011;
		sqrt_table[ 369] = 36'b010011111100111100111000110000110001;
		sqrt_table[ 370] = 36'b010100000000000000000000110000110000;
		sqrt_table[ 371] = 36'b010100000011000011000000110000101110;
		sqrt_table[ 372] = 36'b010100000110000101111000110000101100;
		sqrt_table[ 373] = 36'b010100001001001000101100110000101010;
		sqrt_table[ 374] = 36'b010100001100001011010100110000101001;
		sqrt_table[ 375] = 36'b010100001111001101111000110000100111;
		sqrt_table[ 376] = 36'b010100010010010000010100110000100101;
		sqrt_table[ 377] = 36'b010100010101010010101000110000100011;
		sqrt_table[ 378] = 36'b010100011000010100111000110000100010;
		sqrt_table[ 379] = 36'b010100011011010111000000110000100000;
		sqrt_table[ 380] = 36'b010100011110011001000000110000011110;
		sqrt_table[ 381] = 36'b010100100001011010111000110000011100;
		sqrt_table[ 382] = 36'b010100100100011100101010110000011011;
		sqrt_table[ 383] = 36'b010100100111011110010110110000011001;
		sqrt_table[ 384] = 36'b010100101010011111111000110000010111;
		sqrt_table[ 385] = 36'b010100101101100001011000110000010110;
		sqrt_table[ 386] = 36'b010100110000100010110000110000010011;
		sqrt_table[ 387] = 36'b010100110011100100000000110000010010;
		sqrt_table[ 388] = 36'b010100110110100101001000110000010000;
		sqrt_table[ 389] = 36'b010100111001100110001010110000001111;
		sqrt_table[ 390] = 36'b010100111100100111000110110000001101;
		sqrt_table[ 391] = 36'b010100111111100111111000110000001011;
		sqrt_table[ 392] = 36'b010101000010101000101000110000001001;
		sqrt_table[ 393] = 36'b010101000101101001010000110000001000;
		sqrt_table[ 394] = 36'b010101001000101001110000110000000110;
		sqrt_table[ 395] = 36'b010101001011101010001000110000000100;
		sqrt_table[ 396] = 36'b010101001110101010011010110000000011;
		sqrt_table[ 397] = 36'b010101010001101010100110110000000001;
		sqrt_table[ 398] = 36'b010101010100101010101000101111111111;
		sqrt_table[ 399] = 36'b010101010111101010101000101111111110;
		sqrt_table[ 400] = 36'b010101011010101010100000101111111100;
		sqrt_table[ 401] = 36'b010101011101101010010000101111111010;
		sqrt_table[ 402] = 36'b010101100000101001111010101111111001;
		sqrt_table[ 403] = 36'b010101100011101001011110101111110111;
		sqrt_table[ 404] = 36'b010101100110101000111000101111110101;
		sqrt_table[ 405] = 36'b010101101001101000010000101111110100;
		sqrt_table[ 406] = 36'b010101101100100111100000101111110010;
		sqrt_table[ 407] = 36'b010101101111100110101000101111110000;
		sqrt_table[ 408] = 36'b010101110010100101101100101111101110;
		sqrt_table[ 409] = 36'b010101110101100100100100101111101101;
		sqrt_table[ 410] = 36'b010101111000100011011000101111101011;
		sqrt_table[ 411] = 36'b010101111011100010001000101111101001;
		sqrt_table[ 412] = 36'b010101111110100000110000101111101000;
		sqrt_table[ 413] = 36'b010110000001011111010000101111100110;
		sqrt_table[ 414] = 36'b010110000100011101101010101111100101;
		sqrt_table[ 415] = 36'b010110000111011011111110101111100011;
		sqrt_table[ 416] = 36'b010110001010011010001000101111100001;
		sqrt_table[ 417] = 36'b010110001101011000010000101111100000;
		sqrt_table[ 418] = 36'b010110010000010110010000101111011110;
		sqrt_table[ 419] = 36'b010110010011010100001100101111011100;
		sqrt_table[ 420] = 36'b010110010110010001111100101111011011;
		sqrt_table[ 421] = 36'b010110011001001111101000101111011001;
		sqrt_table[ 422] = 36'b010110011100001101010000101111010111;
		sqrt_table[ 423] = 36'b010110011111001010110000101111010110;
		sqrt_table[ 424] = 36'b010110100010001000001000101111010100;
		sqrt_table[ 425] = 36'b010110100101000101011010101111010011;
		sqrt_table[ 426] = 36'b010110101000000010100110101111010001;
		sqrt_table[ 427] = 36'b010110101010111111101100101111010000;
		sqrt_table[ 428] = 36'b010110101101111100101100101111001110;
		sqrt_table[ 429] = 36'b010110110000111001100100101111001100;
		sqrt_table[ 430] = 36'b010110110011110110010110101111001011;
		sqrt_table[ 431] = 36'b010110110110110011000000101111001001;
		sqrt_table[ 432] = 36'b010110111001101111100100101111000111;
		sqrt_table[ 433] = 36'b010110111100101100000100101111000110;
		sqrt_table[ 434] = 36'b010110111111101000100000101111000100;
		sqrt_table[ 435] = 36'b010111000010100100110000101111000011;
		sqrt_table[ 436] = 36'b010111000101100000111100101111000001;
		sqrt_table[ 437] = 36'b010111001000011101000000101111000000;
		sqrt_table[ 438] = 36'b010111001011011001000000101110111110;
		sqrt_table[ 439] = 36'b010111001110010100111000101110111101;
		sqrt_table[ 440] = 36'b010111010001010000101100101110111011;
		sqrt_table[ 441] = 36'b010111010100001100011000101110111001;
		sqrt_table[ 442] = 36'b010111010111000111111110101110111000;
		sqrt_table[ 443] = 36'b010111011010000011011110101110110110;
		sqrt_table[ 444] = 36'b010111011100111110110110101110110101;
		sqrt_table[ 445] = 36'b010111011111111010001010101110110011;
		sqrt_table[ 446] = 36'b010111100010110101010100101110110001;
		sqrt_table[ 447] = 36'b010111100101110000011100101110110000;
		sqrt_table[ 448] = 36'b010111101000101011100000101110101110;
		sqrt_table[ 449] = 36'b010111101011100110011000101110101101;
		sqrt_table[ 450] = 36'b010111101110100001001100101110101011;
		sqrt_table[ 451] = 36'b010111110001011011111000101110101010;
		sqrt_table[ 452] = 36'b010111110100010110100000101110101000;
		sqrt_table[ 453] = 36'b010111110111010001000100101110100110;
		sqrt_table[ 454] = 36'b010111111010001011011100101110100101;
		sqrt_table[ 455] = 36'b010111111101000101110000101110100011;
		sqrt_table[ 456] = 36'b011000000000000000000000101110100010;
		sqrt_table[ 457] = 36'b011000000010111010001000101110100000;
		sqrt_table[ 458] = 36'b011000000101110100001000101110011111;
		sqrt_table[ 459] = 36'b011000001000101110001000101110011101;
		sqrt_table[ 460] = 36'b011000001011100111111110101110011100;
		sqrt_table[ 461] = 36'b011000001110100001110000101110011010;
		sqrt_table[ 462] = 36'b011000010001011011011000101110011001;
		sqrt_table[ 463] = 36'b011000010100010100111100101110010111;
		sqrt_table[ 464] = 36'b011000010111001110011000101110010110;
		sqrt_table[ 465] = 36'b011000011010000111110000101110010100;
		sqrt_table[ 466] = 36'b011000011101000001000010101110010011;
		sqrt_table[ 467] = 36'b011000011111111010001100101110010001;
		sqrt_table[ 468] = 36'b011000100010110011010100101110001111;
		sqrt_table[ 469] = 36'b011000100101101100010100101110001110;
		sqrt_table[ 470] = 36'b011000101000100101001100101110001101;
		sqrt_table[ 471] = 36'b011000101011011110000000101110001011;
		sqrt_table[ 472] = 36'b011000101110010110101100101110001010;
		sqrt_table[ 473] = 36'b011000110001001111010100101110001000;
		sqrt_table[ 474] = 36'b011000110100000111111000101110000110;
		sqrt_table[ 475] = 36'b011000110111000000010000101110000101;
		sqrt_table[ 476] = 36'b011000111001111000100110101110000100;
		sqrt_table[ 477] = 36'b011000111100110000111000101110000010;
		sqrt_table[ 478] = 36'b011000111111101001000000101110000000;
		sqrt_table[ 479] = 36'b011001000010100001000000101101111111;
		sqrt_table[ 480] = 36'b011001000101011001000000101101111110;
		sqrt_table[ 481] = 36'b011001001000010000111000101101111100;
		sqrt_table[ 482] = 36'b011001001011001000101010101101111011;
		sqrt_table[ 483] = 36'b011001001110000000010100101101111001;
		sqrt_table[ 484] = 36'b011001010000110111111100101101111000;
		sqrt_table[ 485] = 36'b011001010011101111011100101101110110;
		sqrt_table[ 486] = 36'b011001010110100110110110101101110101;
		sqrt_table[ 487] = 36'b011001011001011110001000101101110011;
		sqrt_table[ 488] = 36'b011001011100010101011000101101110010;
		sqrt_table[ 489] = 36'b011001011111001100100000101101110001;
		sqrt_table[ 490] = 36'b011001100010000011100100101101101111;
		sqrt_table[ 491] = 36'b011001100100111010100000101101101110;
		sqrt_table[ 492] = 36'b011001100111110001011000101101101100;
		sqrt_table[ 493] = 36'b011001101010101000001000101101101011;
		sqrt_table[ 494] = 36'b011001101101011110110100101101101001;
		sqrt_table[ 495] = 36'b011001110000010101011000101101100111;
		sqrt_table[ 496] = 36'b011001110011001011111000101101100110;
		sqrt_table[ 497] = 36'b011001110110000010010010101101100101;
		sqrt_table[ 498] = 36'b011001111000111000100110101101100100;
		sqrt_table[ 499] = 36'b011001111011101110110110101101100010;
		sqrt_table[ 500] = 36'b011001111110100101000000101101100000;
		sqrt_table[ 501] = 36'b011010000001011011000000101101011111;
		sqrt_table[ 502] = 36'b011010000100010000111110101101011110;
		sqrt_table[ 503] = 36'b011010000111000110110110101101011100;
		sqrt_table[ 504] = 36'b011010001001111100100110101101011011;
		sqrt_table[ 505] = 36'b011010001100110010010000101101011001;
		sqrt_table[ 506] = 36'b011010001111100111111000101101011000;
		sqrt_table[ 507] = 36'b011010010010011101011100101101010110;
		sqrt_table[ 508] = 36'b011010010101010010110100101101010101;
		sqrt_table[ 509] = 36'b011010011000001000001000101101010011;
		sqrt_table[ 510] = 36'b011010011010111101011000101101010010;
		sqrt_table[ 511] = 36'b011010011101110010100010101101010001;
		sqrt_table[ 512] = 36'b011010100000100111101000101101001111;
		sqrt_table[ 513] = 36'b011010100110010001100000101101001100;
		sqrt_table[ 514] = 36'b011010101011111011000000101101001001;
		sqrt_table[ 515] = 36'b011010110001100100001010101101000110;
		sqrt_table[ 516] = 36'b011010110111001100111100101101000011;
		sqrt_table[ 517] = 36'b011010111100110101011100101101000000;
		sqrt_table[ 518] = 36'b011011000010011101100000101100111110;
		sqrt_table[ 519] = 36'b011011001000000101010100101100111011;
		sqrt_table[ 520] = 36'b011011001101101100101110101100111000;
		sqrt_table[ 521] = 36'b011011010011010011110000101100110101;
		sqrt_table[ 522] = 36'b011011011000111010100000101100110011;
		sqrt_table[ 523] = 36'b011011011110100000111000101100110000;
		sqrt_table[ 524] = 36'b011011100100000110111010101100101101;
		sqrt_table[ 525] = 36'b011011101001101100101000101100101011;
		sqrt_table[ 526] = 36'b011011101111010010000000101100101000;
		sqrt_table[ 527] = 36'b011011110100110111000000101100100101;
		sqrt_table[ 528] = 36'b011011111010011011101100101100100010;
		sqrt_table[ 529] = 36'b011100000000000000000000101100100000;
		sqrt_table[ 530] = 36'b011100000101100100000010101100011101;
		sqrt_table[ 531] = 36'b011100001011000111101110101100011010;
		sqrt_table[ 532] = 36'b011100010000101011000010101100011000;
		sqrt_table[ 533] = 36'b011100010110001110000010101100010101;
		sqrt_table[ 534] = 36'b011100011011110000101100101100010010;
		sqrt_table[ 535] = 36'b011100100001010011000100101100010000;
		sqrt_table[ 536] = 36'b011100100110110101000100101100001101;
		sqrt_table[ 537] = 36'b011100101100010110101100101100001010;
		sqrt_table[ 538] = 36'b011100110001111000000100101100001000;
		sqrt_table[ 539] = 36'b011100110111011001000110101100000101;
		sqrt_table[ 540] = 36'b011100111100111001110000101100000011;
		sqrt_table[ 541] = 36'b011101000010011010001000101100000000;
		sqrt_table[ 542] = 36'b011101000111111010001100101011111101;
		sqrt_table[ 543] = 36'b011101001101011001111000101011111011;
		sqrt_table[ 544] = 36'b011101010010111001010000101011111000;
		sqrt_table[ 545] = 36'b011101011000011000011000101011110101;
		sqrt_table[ 546] = 36'b011101011101110111000110101011110011;
		sqrt_table[ 547] = 36'b011101100011010101100000101011110000;
		sqrt_table[ 548] = 36'b011101101000110011100110101011101110;
		sqrt_table[ 549] = 36'b011101101110010001011010101011101011;
		sqrt_table[ 550] = 36'b011101110011101110111000101011101001;
		sqrt_table[ 551] = 36'b011101111001001100000000101011100110;
		sqrt_table[ 552] = 36'b011101111110101000111000101011100100;
		sqrt_table[ 553] = 36'b011110000100000101011000101011100001;
		sqrt_table[ 554] = 36'b011110001001100001100100101011011111;
		sqrt_table[ 555] = 36'b011110001110111101011100101011011100;
		sqrt_table[ 556] = 36'b011110010100011001000100101011011010;
		sqrt_table[ 557] = 36'b011110011001110100010100101011010111;
		sqrt_table[ 558] = 36'b011110011111001111010000101011010101;
		sqrt_table[ 559] = 36'b011110100100101001111000101011010010;
		sqrt_table[ 560] = 36'b011110101010000100010000101011010000;
		sqrt_table[ 561] = 36'b011110101111011110010000101011001101;
		sqrt_table[ 562] = 36'b011110110100110111111100101011001011;
		sqrt_table[ 563] = 36'b011110111010010001011000101011001000;
		sqrt_table[ 564] = 36'b011110111111101010011100101011000110;
		sqrt_table[ 565] = 36'b011111000101000011010000101011000100;
		sqrt_table[ 566] = 36'b011111001010011011101110101011000001;
		sqrt_table[ 567] = 36'b011111001111110011111100101010111111;
		sqrt_table[ 568] = 36'b011111010101001011110100101010111100;
		sqrt_table[ 569] = 36'b011111011010100011011000101010111010;
		sqrt_table[ 570] = 36'b011111011111111010101000101010111000;
		sqrt_table[ 571] = 36'b011111100101010001101000101010110101;
		sqrt_table[ 572] = 36'b011111101010101000010100101010110011;
		sqrt_table[ 573] = 36'b011111101111111110101100101010110000;
		sqrt_table[ 574] = 36'b011111110101010100110000101010101110;
		sqrt_table[ 575] = 36'b011111111010101010100000101010101011;
		sqrt_table[ 576] = 36'b100000000000000000000010101010101001;
		sqrt_table[ 577] = 36'b100000000101010101001100101010100111;
		sqrt_table[ 578] = 36'b100000001010101010000100101010100100;
		sqrt_table[ 579] = 36'b100000001111111110101010101010100010;
		sqrt_table[ 580] = 36'b100000010101010011000000101010100000;
		sqrt_table[ 581] = 36'b100000011010100111000000101010011101;
		sqrt_table[ 582] = 36'b100000011111111010101110101010011011;
		sqrt_table[ 583] = 36'b100000100101001110001000101010011001;
		sqrt_table[ 584] = 36'b100000101010100001010000101010010110;
		sqrt_table[ 585] = 36'b100000101111110100000110101010010100;
		sqrt_table[ 586] = 36'b100000110101000110101100101010010010;
		sqrt_table[ 587] = 36'b100000111010011000111100101010001111;
		sqrt_table[ 588] = 36'b100000111111101010111010101010001101;
		sqrt_table[ 589] = 36'b100001000100111100100100101010001011;
		sqrt_table[ 590] = 36'b100001001010001110000000101010001001;
		sqrt_table[ 591] = 36'b100001001111011111000100101010000110;
		sqrt_table[ 592] = 36'b100001010100101111111100101010000100;
		sqrt_table[ 593] = 36'b100001011010000000100000101010000010;
		sqrt_table[ 594] = 36'b100001011111010000110000101001111111;
		sqrt_table[ 595] = 36'b100001100100100000101110101001111101;
		sqrt_table[ 596] = 36'b100001101001110000011010101001111011;
		sqrt_table[ 597] = 36'b100001101110111111111000101001111001;
		sqrt_table[ 598] = 36'b100001110100001111000000101001110110;
		sqrt_table[ 599] = 36'b100001111001011101110100101001110100;
		sqrt_table[ 600] = 36'b100001111110101100011100101001110010;
		sqrt_table[ 601] = 36'b100010000011111010101100101001110000;
		sqrt_table[ 602] = 36'b100010001001001000110000101001101110;
		sqrt_table[ 603] = 36'b100010001110010110011100101001101011;
		sqrt_table[ 604] = 36'b100010010011100011111110101001101001;
		sqrt_table[ 605] = 36'b100010011000110001001000101001100111;
		sqrt_table[ 606] = 36'b100010011101111110000100101001100101;
		sqrt_table[ 607] = 36'b100010100011001010101100101001100011;
		sqrt_table[ 608] = 36'b100010101000010111000100101001100000;
		sqrt_table[ 609] = 36'b100010101101100011001010101001011110;
		sqrt_table[ 610] = 36'b100010110010101110111110101001011100;
		sqrt_table[ 611] = 36'b100010110111111010100000101001011010;
		sqrt_table[ 612] = 36'b100010111101000101110100101001011000;
		sqrt_table[ 613] = 36'b100011000010010000110100101001010110;
		sqrt_table[ 614] = 36'b100011000111011011100000101001010011;
		sqrt_table[ 615] = 36'b100011001100100110000010101001010001;
		sqrt_table[ 616] = 36'b100011010001110000001110101001001111;
		sqrt_table[ 617] = 36'b100011010110111010001000101001001101;
		sqrt_table[ 618] = 36'b100011011100000011110100101001001011;
		sqrt_table[ 619] = 36'b100011100001001101001100101001001001;
		sqrt_table[ 620] = 36'b100011100110010110010100101001000111;
		sqrt_table[ 621] = 36'b100011101011011111001100101001000100;
		sqrt_table[ 622] = 36'b100011110000100111110000101001000010;
		sqrt_table[ 623] = 36'b100011110101110000001010101001000000;
		sqrt_table[ 624] = 36'b100011111010111000001110101000111110;
		sqrt_table[ 625] = 36'b100100000000000000000010101000111100;
		sqrt_table[ 626] = 36'b100100000101000111100100101000111010;
		sqrt_table[ 627] = 36'b100100001010001110111000101000111000;
		sqrt_table[ 628] = 36'b100100001111010101111000101000110110;
		sqrt_table[ 629] = 36'b100100010100011100101000101000110100;
		sqrt_table[ 630] = 36'b100100011001100011001000101000110010;
		sqrt_table[ 631] = 36'b100100011110101001011000101000110000;
		sqrt_table[ 632] = 36'b100100100011101111011000101000101101;
		sqrt_table[ 633] = 36'b100100101000110101001000101000101100;
		sqrt_table[ 634] = 36'b100100101101111010100110101000101001;
		sqrt_table[ 635] = 36'b100100110010111111110100101000100111;
		sqrt_table[ 636] = 36'b100100111000000100110000101000100101;
		sqrt_table[ 637] = 36'b100100111101001001011110101000100011;
		sqrt_table[ 638] = 36'b100101000010001101111000101000100001;
		sqrt_table[ 639] = 36'b100101000111010010001010101000011111;
		sqrt_table[ 640] = 36'b100101001100010110000110101000011101;
		sqrt_table[ 641] = 36'b100101010001011001110010101000011011;
		sqrt_table[ 642] = 36'b100101010110011101001110101000011001;
		sqrt_table[ 643] = 36'b100101011011100000011010101000010111;
		sqrt_table[ 644] = 36'b100101100000100011010110101000010101;
		sqrt_table[ 645] = 36'b100101100101100110000010101000010011;
		sqrt_table[ 646] = 36'b100101101010101000011110101000010001;
		sqrt_table[ 647] = 36'b100101101111101010101010101000001111;
		sqrt_table[ 648] = 36'b100101110100101100100110101000001101;
		sqrt_table[ 649] = 36'b100101111001101110010010101000001011;
		sqrt_table[ 650] = 36'b100101111110101111101110101000001001;
		sqrt_table[ 651] = 36'b100110000011110000111010101000000111;
		sqrt_table[ 652] = 36'b100110001000110001110100101000000101;
		sqrt_table[ 653] = 36'b100110001101110010100010101000000011;
		sqrt_table[ 654] = 36'b100110010010110011000000101000000001;
		sqrt_table[ 655] = 36'b100110010111110011001100100111111111;
		sqrt_table[ 656] = 36'b100110011100110011001000100111111101;
		sqrt_table[ 657] = 36'b100110100001110010111000100111111011;
		sqrt_table[ 658] = 36'b100110100110110010011000100111111010;
		sqrt_table[ 659] = 36'b100110101011110001101000100111111000;
		sqrt_table[ 660] = 36'b100110110000110000101000100111110110;
		sqrt_table[ 661] = 36'b100110110101101111011000100111110100;
		sqrt_table[ 662] = 36'b100110111010101101111000100111110010;
		sqrt_table[ 663] = 36'b100110111111101100001000100111110000;
		sqrt_table[ 664] = 36'b100111000100101010001100100111101110;
		sqrt_table[ 665] = 36'b100111001001100111111110100111101100;
		sqrt_table[ 666] = 36'b100111001110100101100010100111101010;
		sqrt_table[ 667] = 36'b100111010011100010110110100111101000;
		sqrt_table[ 668] = 36'b100111011000011111111000100111100110;
		sqrt_table[ 669] = 36'b100111011101011100110000100111100100;
		sqrt_table[ 670] = 36'b100111100010011001010100100111100011;
		sqrt_table[ 671] = 36'b100111100111010101101100100111100001;
		sqrt_table[ 672] = 36'b100111101100010001110100100111011111;
		sqrt_table[ 673] = 36'b100111110001001101110000100111011101;
		sqrt_table[ 674] = 36'b100111110110001001011010100111011011;
		sqrt_table[ 675] = 36'b100111111011000100110110100111011001;
		sqrt_table[ 676] = 36'b101000000000000000000000100111010111;
		sqrt_table[ 677] = 36'b101000000100111010111100100111010101;
		sqrt_table[ 678] = 36'b101000001001110101101100100111010100;
		sqrt_table[ 679] = 36'b101000001110110000001100100111010010;
		sqrt_table[ 680] = 36'b101000010011101010011100100111010000;
		sqrt_table[ 681] = 36'b101000011000100100011110100111001110;
		sqrt_table[ 682] = 36'b101000011101011110010010100111001100;
		sqrt_table[ 683] = 36'b101000100010010111111000100111001010;
		sqrt_table[ 684] = 36'b101000100111010001001100100111001001;
		sqrt_table[ 685] = 36'b101000101100001010010100100111000111;
		sqrt_table[ 686] = 36'b101000110001000011001110100111000101;
		sqrt_table[ 687] = 36'b101000110101111011111000100111000011;
		sqrt_table[ 688] = 36'b101000111010110100010000100111000001;
		sqrt_table[ 689] = 36'b101000111111101100100000100110111111;
		sqrt_table[ 690] = 36'b101001000100100100100000100110111110;
		sqrt_table[ 691] = 36'b101001001001011100010000100110111100;
		sqrt_table[ 692] = 36'b101001001110010011110010100110111010;
		sqrt_table[ 693] = 36'b101001010011001011000110100110111000;
		sqrt_table[ 694] = 36'b101001011000000010001000100110110110;
		sqrt_table[ 695] = 36'b101001011100111001000000100110110101;
		sqrt_table[ 696] = 36'b101001100001101111101000100110110011;
		sqrt_table[ 697] = 36'b101001100110100110000010100110110001;
		sqrt_table[ 698] = 36'b101001101011011100001100100110101111;
		sqrt_table[ 699] = 36'b101001110000010010001100100110101110;
		sqrt_table[ 700] = 36'b101001110101000111111100100110101100;
		sqrt_table[ 701] = 36'b101001111001111101011010100110101010;
		sqrt_table[ 702] = 36'b101001111110110010101110100110101000;
		sqrt_table[ 703] = 36'b101010000011100111110100100110100111;
		sqrt_table[ 704] = 36'b101010001000011100101100100110100101;
		sqrt_table[ 705] = 36'b101010001101010001010100100110100011;
		sqrt_table[ 706] = 36'b101010010010000101101100100110100001;
		sqrt_table[ 707] = 36'b101010010110111001111000100110011111;
		sqrt_table[ 708] = 36'b101010011011101101111000100110011110;
		sqrt_table[ 709] = 36'b101010100000100001101100100110011100;
		sqrt_table[ 710] = 36'b101010100101010101001100100110011010;
		sqrt_table[ 711] = 36'b101010101010001000100100100110011001;
		sqrt_table[ 712] = 36'b101010101110111011101100100110010111;
		sqrt_table[ 713] = 36'b101010110011101110100100100110010101;
		sqrt_table[ 714] = 36'b101010111000100001010000100110010100;
		sqrt_table[ 715] = 36'b101010111101010011110000100110010010;
		sqrt_table[ 716] = 36'b101011000010000110000000100110010000;
		sqrt_table[ 717] = 36'b101011000110111000000000100110001110;
		sqrt_table[ 718] = 36'b101011001011101001110100100110001100;
		sqrt_table[ 719] = 36'b101011010000011011011100100110001011;
		sqrt_table[ 720] = 36'b101011010101001100110110100110001001;
		sqrt_table[ 721] = 36'b101011011001111110000100100110001000;
		sqrt_table[ 722] = 36'b101011011110101111000100100110000110;
		sqrt_table[ 723] = 36'b101011100011011111110010100110000100;
		sqrt_table[ 724] = 36'b101011101000010000011000100110000010;
		sqrt_table[ 725] = 36'b101011101101000000101100100110000001;
		sqrt_table[ 726] = 36'b101011110001110000110110100101111111;
		sqrt_table[ 727] = 36'b101011110110100000110000100101111101;
		sqrt_table[ 728] = 36'b101011111011010000100000100101111100;
		sqrt_table[ 729] = 36'b101100000000000000000010100101111010;
		sqrt_table[ 730] = 36'b101100000100101111010100100101111000;
		sqrt_table[ 731] = 36'b101100001001011110011100100101110111;
		sqrt_table[ 732] = 36'b101100001110001101010010100101110101;
		sqrt_table[ 733] = 36'b101100010010111011111100100101110011;
		sqrt_table[ 734] = 36'b101100010111101010011100100101110010;
		sqrt_table[ 735] = 36'b101100011100011000101110100101110000;
		sqrt_table[ 736] = 36'b101100100001000110110000100101101110;
		sqrt_table[ 737] = 36'b101100100101110100101000100101101101;
		sqrt_table[ 738] = 36'b101100101010100010010000100101101011;
		sqrt_table[ 739] = 36'b101100101111001111110000100101101010;
		sqrt_table[ 740] = 36'b101100110011111101000000100101101000;
		sqrt_table[ 741] = 36'b101100111000101010000000100101100110;
		sqrt_table[ 742] = 36'b101100111101010110111000100101100101;
		sqrt_table[ 743] = 36'b101101000010000011100010100101100011;
		sqrt_table[ 744] = 36'b101101000110101111111100100101100001;
		sqrt_table[ 745] = 36'b101101001011011100001100100101100000;
		sqrt_table[ 746] = 36'b101101010000001000001100100101011110;
		sqrt_table[ 747] = 36'b101101010100110100000100100101011101;
		sqrt_table[ 748] = 36'b101101011001011111101010100101011011;
		sqrt_table[ 749] = 36'b101101011110001011000100100101011001;
		sqrt_table[ 750] = 36'b101101100010110110010100100101011000;
		sqrt_table[ 751] = 36'b101101100111100001010100100101010110;
		sqrt_table[ 752] = 36'b101101101100001100001100100101010101;
		sqrt_table[ 753] = 36'b101101110000110110110110100101010011;
		sqrt_table[ 754] = 36'b101101110101100001010000100101010001;
		sqrt_table[ 755] = 36'b101101111010001011011110100101010000;
		sqrt_table[ 756] = 36'b101101111110110101100000100101001110;
		sqrt_table[ 757] = 36'b101110000011011111011000100101001101;
		sqrt_table[ 758] = 36'b101110001000001001000000100101001011;
		sqrt_table[ 759] = 36'b101110001100110010011110100101001010;
		sqrt_table[ 760] = 36'b101110010001011011101110100101001000;
		sqrt_table[ 761] = 36'b101110010110000100110000100101000110;
		sqrt_table[ 762] = 36'b101110011010101101101000100101000101;
		sqrt_table[ 763] = 36'b101110011111010110010100100101000100;
		sqrt_table[ 764] = 36'b101110100011111110110100100101000010;
		sqrt_table[ 765] = 36'b101110101000100111000110100101000000;
		sqrt_table[ 766] = 36'b101110101101001111001000100100111111;
		sqrt_table[ 767] = 36'b101110110001110111000010100100111101;
		sqrt_table[ 768] = 36'b101110110110011110110000100100111100;
		sqrt_table[ 769] = 36'b101110111011000110001100100100111010;
		sqrt_table[ 770] = 36'b101110111111101101100100100100111001;
		sqrt_table[ 771] = 36'b101111000100010100101100100100110111;
		sqrt_table[ 772] = 36'b101111001000111011101000100100110110;
		sqrt_table[ 773] = 36'b101111001101100010010110100100110100;
		sqrt_table[ 774] = 36'b101111010010001000111000100100110010;
		sqrt_table[ 775] = 36'b101111010110101111010010100100110001;
		sqrt_table[ 776] = 36'b101111011011010101011100100100101111;
		sqrt_table[ 777] = 36'b101111011111111011011100100100101110;
		sqrt_table[ 778] = 36'b101111100100100001001100100100101101;
		sqrt_table[ 779] = 36'b101111101001000110110100100100101011;
		sqrt_table[ 780] = 36'b101111101101101100001100100100101001;
		sqrt_table[ 781] = 36'b101111110010010001011100100100101000;
		sqrt_table[ 782] = 36'b101111110110110110100000100100100111;
		sqrt_table[ 783] = 36'b101111111011011011011000100100100101;
		sqrt_table[ 784] = 36'b110000000000000000000000100100100011;
		sqrt_table[ 785] = 36'b110000000100100100011110100100100010;
		sqrt_table[ 786] = 36'b110000001001001000110000100100100000;
		sqrt_table[ 787] = 36'b110000001101101100111000100100011111;
		sqrt_table[ 788] = 36'b110000010010010000110100100100011110;
		sqrt_table[ 789] = 36'b110000010110110100100010100100011100;
		sqrt_table[ 790] = 36'b110000011011011000000100100100011010;
		sqrt_table[ 791] = 36'b110000011111111011011110100100011001;
		sqrt_table[ 792] = 36'b110000100100011110101000100100011000;
		sqrt_table[ 793] = 36'b110000101001000001101010100100010110;
		sqrt_table[ 794] = 36'b110000101101100100011100100100010101;
		sqrt_table[ 795] = 36'b110000110010000111000100100100010011;
		sqrt_table[ 796] = 36'b110000110110101001100100100100010010;
		sqrt_table[ 797] = 36'b110000111011001011110000100100010000;
		sqrt_table[ 798] = 36'b110000111111101101111000100100001111;
		sqrt_table[ 799] = 36'b110001000100001111110000100100001101;
		sqrt_table[ 800] = 36'b110001001000110001100000100100001100;
		sqrt_table[ 801] = 36'b110001001101010011000100100100001011;
		sqrt_table[ 802] = 36'b110001010001110100011010100100001001;
		sqrt_table[ 803] = 36'b110001010110010101100110100100001000;
		sqrt_table[ 804] = 36'b110001011010110110100110100100000110;
		sqrt_table[ 805] = 36'b110001011111010111011100100100000101;
		sqrt_table[ 806] = 36'b110001100011111000000000100100000011;
		sqrt_table[ 807] = 36'b110001101000011000100000100100000010;
		sqrt_table[ 808] = 36'b110001101100111000110000100100000000;
		sqrt_table[ 809] = 36'b110001110001011000111010100011111111;
		sqrt_table[ 810] = 36'b110001110101111000110100100011111110;
		sqrt_table[ 811] = 36'b110001111010011000100110100011111100;
		sqrt_table[ 812] = 36'b110001111110111000001000100011111011;
		sqrt_table[ 813] = 36'b110010000011010111100000100011111001;
		sqrt_table[ 814] = 36'b110010000111110110110000100011111000;
		sqrt_table[ 815] = 36'b110010001100010101110100100011110111;
		sqrt_table[ 816] = 36'b110010010000110100101010100011110101;
		sqrt_table[ 817] = 36'b110010010101010011011000100011110100;
		sqrt_table[ 818] = 36'b110010011001110001111000100011110010;
		sqrt_table[ 819] = 36'b110010011110010000001110100011110001;
		sqrt_table[ 820] = 36'b110010100010101110011000100011101111;
		sqrt_table[ 821] = 36'b110010100111001100010110100011101110;
		sqrt_table[ 822] = 36'b110010101011101010001100100011101101;
		sqrt_table[ 823] = 36'b110010110000000111110100100011101011;
		sqrt_table[ 824] = 36'b110010110100100101010100100011101010;
		sqrt_table[ 825] = 36'b110010111001000010100100100011101001;
		sqrt_table[ 826] = 36'b110010111101011111101100100011100111;
		sqrt_table[ 827] = 36'b110011000001111100101100100011100110;
		sqrt_table[ 828] = 36'b110011000110011001011100100011100100;
		sqrt_table[ 829] = 36'b110011001010110110000010100011100011;
		sqrt_table[ 830] = 36'b110011001111010010100000100011100010;
		sqrt_table[ 831] = 36'b110011010011101110101100100011100000;
		sqrt_table[ 832] = 36'b110011011000001010110110100011011111;
		sqrt_table[ 833] = 36'b110011011100100110110000100011011110;
		sqrt_table[ 834] = 36'b110011100001000010100010100011011100;
		sqrt_table[ 835] = 36'b110011100101011110000100100011011011;
		sqrt_table[ 836] = 36'b110011101001111001100000100011011010;
		sqrt_table[ 837] = 36'b110011101110010100101110100011011000;
		sqrt_table[ 838] = 36'b110011110010101111110100100011010111;
		sqrt_table[ 839] = 36'b110011110111001010101100100011010110;
		sqrt_table[ 840] = 36'b110011111011100101011110100011010100;
		sqrt_table[ 841] = 36'b110100000000000000000000100011010011;
		sqrt_table[ 842] = 36'b110100000100011010011000100011010001;
		sqrt_table[ 843] = 36'b110100001000110100101010100011010000;
		sqrt_table[ 844] = 36'b110100001101001110101100100011001111;
		sqrt_table[ 845] = 36'b110100010001101000100100100011001101;
		sqrt_table[ 846] = 36'b110100010110000010010110100011001100;
		sqrt_table[ 847] = 36'b110100011010011011111000100011001011;
		sqrt_table[ 848] = 36'b110100011110110101010000100011001001;
		sqrt_table[ 849] = 36'b110100100011001110100000100011001000;
		sqrt_table[ 850] = 36'b110100100111100111101000100011000111;
		sqrt_table[ 851] = 36'b110100101100000000100000100011000110;
		sqrt_table[ 852] = 36'b110100110000011001001110100011000100;
		sqrt_table[ 853] = 36'b110100110100110001110100100011000011;
		sqrt_table[ 854] = 36'b110100111001001010001100100011000010;
		sqrt_table[ 855] = 36'b110100111101100010011110100011000000;
		sqrt_table[ 856] = 36'b110101000001111010100010100010111111;
		sqrt_table[ 857] = 36'b110101000110010010011100100010111110;
		sqrt_table[ 858] = 36'b110101001010101010001100100010111100;
		sqrt_table[ 859] = 36'b110101001111000001110100100010111011;
		sqrt_table[ 860] = 36'b110101010011011001001100100010111010;
		sqrt_table[ 861] = 36'b110101010111110000011100100010111000;
		sqrt_table[ 862] = 36'b110101011100000111100110100010110111;
		sqrt_table[ 863] = 36'b110101100000011110100000100010110110;
		sqrt_table[ 864] = 36'b110101100100110101010010100010110101;
		sqrt_table[ 865] = 36'b110101101001001011111010100010110011;
		sqrt_table[ 866] = 36'b110101101101100010010110100010110010;
		sqrt_table[ 867] = 36'b110101110001111000101100100010110001;
		sqrt_table[ 868] = 36'b110101110110001110110000100010101111;
		sqrt_table[ 869] = 36'b110101111010100100110010100010101110;
		sqrt_table[ 870] = 36'b110101111110111010100100100010101101;
		sqrt_table[ 871] = 36'b110110000011010000010000100010101100;
		sqrt_table[ 872] = 36'b110110000111100101101100100010101010;
		sqrt_table[ 873] = 36'b110110001011111011000100100010101001;
		sqrt_table[ 874] = 36'b110110010000010000010000100010101000;
		sqrt_table[ 875] = 36'b110110010100100101010000100010100111;
		sqrt_table[ 876] = 36'b110110011000111010001010100010100101;
		sqrt_table[ 877] = 36'b110110011101001110110110100010100100;
		sqrt_table[ 878] = 36'b110110100001100011011000100010100011;
		sqrt_table[ 879] = 36'b110110100101110111110000100010100001;
		sqrt_table[ 880] = 36'b110110101010001011111100100010100000;
		sqrt_table[ 881] = 36'b110110101110100000000100100010011111;
		sqrt_table[ 882] = 36'b110110110010110100000000100010011110;
		sqrt_table[ 883] = 36'b110110110111000111110000100010011100;
		sqrt_table[ 884] = 36'b110110111011011011010110100010011011;
		sqrt_table[ 885] = 36'b110110111111101110110010100010011010;
		sqrt_table[ 886] = 36'b110111000100000010000110100010011001;
		sqrt_table[ 887] = 36'b110111001000010101001110100010011000;
		sqrt_table[ 888] = 36'b110111001100101000001110100010010110;
		sqrt_table[ 889] = 36'b110111010000111011000010100010010101;
		sqrt_table[ 890] = 36'b110111010101001101110000100010010100;
		sqrt_table[ 891] = 36'b110111011001100000010000100010010011;
		sqrt_table[ 892] = 36'b110111011101110010100100100010010001;
		sqrt_table[ 893] = 36'b110111100010000100110100100010010000;
		sqrt_table[ 894] = 36'b110111100110010110111000100010001111;
		sqrt_table[ 895] = 36'b110111101010101000110000100010001110;
		sqrt_table[ 896] = 36'b110111101110111010100000100010001100;
		sqrt_table[ 897] = 36'b110111110011001100001000100010001011;
		sqrt_table[ 898] = 36'b110111110111011101100100100010001010;
		sqrt_table[ 899] = 36'b110111111011101110111000100010001001;
		sqrt_table[ 900] = 36'b111000000000000000000000100010001000;
		sqrt_table[ 901] = 36'b111000000100010001000000100010000110;
		sqrt_table[ 902] = 36'b111000001000100001110110100010000101;
		sqrt_table[ 903] = 36'b111000001100110010100100100010000100;
		sqrt_table[ 904] = 36'b111000010001000011000100100010000011;
		sqrt_table[ 905] = 36'b111000010101010011011100100010000010;
		sqrt_table[ 906] = 36'b111000011001100011101110100010000000;
		sqrt_table[ 907] = 36'b111000011101110011110010100001111111;
		sqrt_table[ 908] = 36'b111000100010000011101110100001111110;
		sqrt_table[ 909] = 36'b111000100110010011100000100001111101;
		sqrt_table[ 910] = 36'b111000101010100011001000100001111100;
		sqrt_table[ 911] = 36'b111000101110110010101010100001111010;
		sqrt_table[ 912] = 36'b111000110011000001111110100001111001;
		sqrt_table[ 913] = 36'b111000110111010001001010100001111000;
		sqrt_table[ 914] = 36'b111000111011100000001100100001110111;
		sqrt_table[ 915] = 36'b111000111111101111000100100001110110;
		sqrt_table[ 916] = 36'b111001000011111101110100100001110100;
		sqrt_table[ 917] = 36'b111001001000001100011000100001110011;
		sqrt_table[ 918] = 36'b111001001100011010111000100001110010;
		sqrt_table[ 919] = 36'b111001010000101001001100100001110001;
		sqrt_table[ 920] = 36'b111001010100110111010100100001110000;
		sqrt_table[ 921] = 36'b111001011001000101010100100001101110;
		sqrt_table[ 922] = 36'b111001011101010011001100100001101101;
		sqrt_table[ 923] = 36'b111001100001100000111010100001101100;
		sqrt_table[ 924] = 36'b111001100101101110011110100001101011;
		sqrt_table[ 925] = 36'b111001101001111011111100100001101010;
		sqrt_table[ 926] = 36'b111001101110001001001100100001101001;
		sqrt_table[ 927] = 36'b111001110010010110010100100001101000;
		sqrt_table[ 928] = 36'b111001110110100011010100100001100110;
		sqrt_table[ 929] = 36'b111001111010110000001010100001100101;
		sqrt_table[ 930] = 36'b111001111110111100110110100001100100;
		sqrt_table[ 931] = 36'b111010000011001001011100100001100011;
		sqrt_table[ 932] = 36'b111010000111010101110100100001100010;
		sqrt_table[ 933] = 36'b111010001011100010000100100001100001;
		sqrt_table[ 934] = 36'b111010001111101110001100100001100000;
		sqrt_table[ 935] = 36'b111010010011111010001110100001011110;
		sqrt_table[ 936] = 36'b111010011000000110000000100001011101;
		sqrt_table[ 937] = 36'b111010011100010001110000100001011100;
		sqrt_table[ 938] = 36'b111010100000011101010000100001011011;
		sqrt_table[ 939] = 36'b111010100100101000101100100001011010;
		sqrt_table[ 940] = 36'b111010101000110011111100100001011001;
		sqrt_table[ 941] = 36'b111010101100111111000100100001010111;
		sqrt_table[ 942] = 36'b111010110001001010000000100001010110;
		sqrt_table[ 943] = 36'b111010110101010100111010100001010101;
		sqrt_table[ 944] = 36'b111010111001011111100110100001010100;
		sqrt_table[ 945] = 36'b111010111101101010001000100001010011;
		sqrt_table[ 946] = 36'b111011000001110100100100100001010010;
		sqrt_table[ 947] = 36'b111011000101111110110100100001010001;
		sqrt_table[ 948] = 36'b111011001010001000111100100001010000;
		sqrt_table[ 949] = 36'b111011001110010010111100100001001110;
		sqrt_table[ 950] = 36'b111011010010011100110000100001001101;
		sqrt_table[ 951] = 36'b111011010110100110100000100001001100;
		sqrt_table[ 952] = 36'b111011011010110000000110100001001011;
		sqrt_table[ 953] = 36'b111011011110111001100100100001001010;
		sqrt_table[ 954] = 36'b111011100011000010110100100001001001;
		sqrt_table[ 955] = 36'b111011100111001100000000100001001000;
		sqrt_table[ 956] = 36'b111011101011010101000000100001000111;
		sqrt_table[ 957] = 36'b111011101111011101111000100001000101;
		sqrt_table[ 958] = 36'b111011110011100110101000100001000101;
		sqrt_table[ 959] = 36'b111011110111101111001100100001000011;
		sqrt_table[ 960] = 36'b111011111011110111101100100001000010;
		sqrt_table[ 961] = 36'b111100000000000000000010100001000001;
		sqrt_table[ 962] = 36'b111100000100001000001100100001000000;
		sqrt_table[ 963] = 36'b111100001000010000010000100000111111;
		sqrt_table[ 964] = 36'b111100001100011000001100100000111110;
		sqrt_table[ 965] = 36'b111100010000011111111100100000111101;
		sqrt_table[ 966] = 36'b111100010100100111100100100000111100;
		sqrt_table[ 967] = 36'b111100011000101111000100100000111010;
		sqrt_table[ 968] = 36'b111100011100110110011100100000111010;
		sqrt_table[ 969] = 36'b111100100000111101101100100000111000;
		sqrt_table[ 970] = 36'b111100100101000100110000100000110111;
		sqrt_table[ 971] = 36'b111100101001001011110000100000110110;
		sqrt_table[ 972] = 36'b111100101101010010100110100000110101;
		sqrt_table[ 973] = 36'b111100110001011001010010100000110100;
		sqrt_table[ 974] = 36'b111100110101011111110100100000110011;
		sqrt_table[ 975] = 36'b111100111001100110010000100000110010;
		sqrt_table[ 976] = 36'b111100111101101100100100100000110001;
		sqrt_table[ 977] = 36'b111101000001110010101100100000110000;
		sqrt_table[ 978] = 36'b111101000101111000101100100000101111;
		sqrt_table[ 979] = 36'b111101001001111110100100100000101110;
		sqrt_table[ 980] = 36'b111101001110000100010100100000101100;
		sqrt_table[ 981] = 36'b111101010010001001111100100000101100;
		sqrt_table[ 982] = 36'b111101010110001111011100100000101010;
		sqrt_table[ 983] = 36'b111101011010010100110000100000101001;
		sqrt_table[ 984] = 36'b111101011110011010000000100000101000;
		sqrt_table[ 985] = 36'b111101100010011111000110100000100111;
		sqrt_table[ 986] = 36'b111101100110100100000010100000100110;
		sqrt_table[ 987] = 36'b111101101010101000110110100000100101;
		sqrt_table[ 988] = 36'b111101101110101101100010100000100100;
		sqrt_table[ 989] = 36'b111101110010110010000110100000100011;
		sqrt_table[ 990] = 36'b111101110110110110100100100000100010;
		sqrt_table[ 991] = 36'b111101111010111010110100100000100001;
		sqrt_table[ 992] = 36'b111101111110111111000000100000100000;
		sqrt_table[ 993] = 36'b111110000011000011000000100000011111;
		sqrt_table[ 994] = 36'b111110000111000110111100100000011110;
		sqrt_table[ 995] = 36'b111110001011001010101100100000011101;
		sqrt_table[ 996] = 36'b111110001111001110010100100000011100;
		sqrt_table[ 997] = 36'b111110010011010001110100100000011011;
		sqrt_table[ 998] = 36'b111110010111010101001110100000011010;
		sqrt_table[ 999] = 36'b111110011011011000011100100000011000;
		sqrt_table[1000] = 36'b111110011111011011100100100000011000;
		sqrt_table[1001] = 36'b111110100011011110100100100000010110;
		sqrt_table[1002] = 36'b111110100111100001011100100000010110;
		sqrt_table[1003] = 36'b111110101011100100001000100000010100;
		sqrt_table[1004] = 36'b111110101111100110110000100000010011;
		sqrt_table[1005] = 36'b111110110011101001001100100000010010;
		sqrt_table[1006] = 36'b111110110111101011100100100000010001;
		sqrt_table[1007] = 36'b111110111011101101110000100000010000;
		sqrt_table[1008] = 36'b111110111111101111111000100000001111;
		sqrt_table[1009] = 36'b111111000011110001110110100000001110;
		sqrt_table[1010] = 36'b111111000111110011101000100000001101;
		sqrt_table[1011] = 36'b111111001011110101011010100000001100;
		sqrt_table[1012] = 36'b111111001111110110111100100000001011;
		sqrt_table[1013] = 36'b111111010011111000011010100000001010;
		sqrt_table[1014] = 36'b111111010111111001101110100000001001;
		sqrt_table[1015] = 36'b111111011011111010111010100000001000;
		sqrt_table[1016] = 36'b111111011111111011111100100000000111;
		sqrt_table[1017] = 36'b111111100011111100111100100000000110;
		sqrt_table[1018] = 36'b111111100111111101110000100000000101;
		sqrt_table[1019] = 36'b111111101011111110011100100000000100;
		sqrt_table[1020] = 36'b111111101111111111000000100000000011;
		sqrt_table[1021] = 36'b111111110011111111011100100000000010;
		sqrt_table[1022] = 36'b111111110111111111110000100000000001;
		sqrt_table[1023] = 36'b111111111011111111111100100000000000;
	end
endmodule

`default_nettype wire